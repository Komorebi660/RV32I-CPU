// Copyright (c) 2022 Komorebi660
// Functional Test file name: ../binary/1testAll.data

module mem #(                    
    parameter  ADDR_LEN  = 11    
) (
    input  clk, rst,
    input  [ADDR_LEN-1:0] addr, // memory address
    output reg [31:0] rd_data,  // data read out
    input  wr_req,              // write request
    input  [31:0] wr_data       // data write in
);
localparam MEM_SIZE = 1<<ADDR_LEN;
reg [31:0] ram_cell [MEM_SIZE];

always @ (posedge clk or posedge rst)
    if(rst)
        rd_data <= 0;
    else
        rd_data <= ram_cell[addr];

always @ (posedge clk)
    if(wr_req) 
        ram_cell[addr] <= wr_data;

initial begin
        ram_cell[       0] = 32'h00000013;
        ram_cell[       1] = 32'h00000093;
        ram_cell[       2] = 32'h00000113;
        ram_cell[       3] = 32'h00208f33;
        ram_cell[       4] = 32'h00000e93;
        ram_cell[       5] = 32'h00200193;
        ram_cell[       6] = 32'h01df0463;
        ram_cell[       7] = 32'h2ac0206f;
        ram_cell[       8] = 32'h00100093;
        ram_cell[       9] = 32'h00100113;
        ram_cell[      10] = 32'h00208f33;
        ram_cell[      11] = 32'h00200e93;
        ram_cell[      12] = 32'h00300193;
        ram_cell[      13] = 32'h01df0463;
        ram_cell[      14] = 32'h2900206f;
        ram_cell[      15] = 32'h00300093;
        ram_cell[      16] = 32'h00700113;
        ram_cell[      17] = 32'h00208f33;
        ram_cell[      18] = 32'h00a00e93;
        ram_cell[      19] = 32'h00400193;
        ram_cell[      20] = 32'h01df0463;
        ram_cell[      21] = 32'h2740206f;
        ram_cell[      22] = 32'h00000093;
        ram_cell[      23] = 32'hffff8137;
        ram_cell[      24] = 32'h00208f33;
        ram_cell[      25] = 32'hffff8eb7;
        ram_cell[      26] = 32'h00500193;
        ram_cell[      27] = 32'h01df0463;
        ram_cell[      28] = 32'h2580206f;
        ram_cell[      29] = 32'h800000b7;
        ram_cell[      30] = 32'h00000113;
        ram_cell[      31] = 32'h00208f33;
        ram_cell[      32] = 32'h80000eb7;
        ram_cell[      33] = 32'h00600193;
        ram_cell[      34] = 32'h01df0463;
        ram_cell[      35] = 32'h23c0206f;
        ram_cell[      36] = 32'h800000b7;
        ram_cell[      37] = 32'hffff8137;
        ram_cell[      38] = 32'h00208f33;
        ram_cell[      39] = 32'h7fff8eb7;
        ram_cell[      40] = 32'h00700193;
        ram_cell[      41] = 32'h01df0463;
        ram_cell[      42] = 32'h2200206f;
        ram_cell[      43] = 32'h00000093;
        ram_cell[      44] = 32'h00008137;
        ram_cell[      45] = 32'hfff10113;
        ram_cell[      46] = 32'h00208f33;
        ram_cell[      47] = 32'h00008eb7;
        ram_cell[      48] = 32'hfffe8e93;
        ram_cell[      49] = 32'h00800193;
        ram_cell[      50] = 32'h01df0463;
        ram_cell[      51] = 32'h1fc0206f;
        ram_cell[      52] = 32'h800000b7;
        ram_cell[      53] = 32'hfff08093;
        ram_cell[      54] = 32'h00000113;
        ram_cell[      55] = 32'h00208f33;
        ram_cell[      56] = 32'h80000eb7;
        ram_cell[      57] = 32'hfffe8e93;
        ram_cell[      58] = 32'h00900193;
        ram_cell[      59] = 32'h01df0463;
        ram_cell[      60] = 32'h1d80206f;
        ram_cell[      61] = 32'h800000b7;
        ram_cell[      62] = 32'hfff08093;
        ram_cell[      63] = 32'h00008137;
        ram_cell[      64] = 32'hfff10113;
        ram_cell[      65] = 32'h00208f33;
        ram_cell[      66] = 32'h80008eb7;
        ram_cell[      67] = 32'hffee8e93;
        ram_cell[      68] = 32'h00a00193;
        ram_cell[      69] = 32'h01df0463;
        ram_cell[      70] = 32'h1b00206f;
        ram_cell[      71] = 32'h800000b7;
        ram_cell[      72] = 32'h00008137;
        ram_cell[      73] = 32'hfff10113;
        ram_cell[      74] = 32'h00208f33;
        ram_cell[      75] = 32'h80008eb7;
        ram_cell[      76] = 32'hfffe8e93;
        ram_cell[      77] = 32'h00b00193;
        ram_cell[      78] = 32'h01df0463;
        ram_cell[      79] = 32'h18c0206f;
        ram_cell[      80] = 32'h800000b7;
        ram_cell[      81] = 32'hfff08093;
        ram_cell[      82] = 32'hffff8137;
        ram_cell[      83] = 32'h00208f33;
        ram_cell[      84] = 32'h7fff8eb7;
        ram_cell[      85] = 32'hfffe8e93;
        ram_cell[      86] = 32'h00c00193;
        ram_cell[      87] = 32'h01df0463;
        ram_cell[      88] = 32'h1680206f;
        ram_cell[      89] = 32'h00000093;
        ram_cell[      90] = 32'hfff00113;
        ram_cell[      91] = 32'h00208f33;
        ram_cell[      92] = 32'hfff00e93;
        ram_cell[      93] = 32'h00d00193;
        ram_cell[      94] = 32'h01df0463;
        ram_cell[      95] = 32'h14c0206f;
        ram_cell[      96] = 32'hfff00093;
        ram_cell[      97] = 32'h00100113;
        ram_cell[      98] = 32'h00208f33;
        ram_cell[      99] = 32'h00000e93;
        ram_cell[     100] = 32'h00e00193;
        ram_cell[     101] = 32'h01df0463;
        ram_cell[     102] = 32'h1300206f;
        ram_cell[     103] = 32'hfff00093;
        ram_cell[     104] = 32'hfff00113;
        ram_cell[     105] = 32'h00208f33;
        ram_cell[     106] = 32'hffe00e93;
        ram_cell[     107] = 32'h00f00193;
        ram_cell[     108] = 32'h01df0463;
        ram_cell[     109] = 32'h1140206f;
        ram_cell[     110] = 32'h00100093;
        ram_cell[     111] = 32'h80000137;
        ram_cell[     112] = 32'hfff10113;
        ram_cell[     113] = 32'h00208f33;
        ram_cell[     114] = 32'h80000eb7;
        ram_cell[     115] = 32'h01000193;
        ram_cell[     116] = 32'h01df0463;
        ram_cell[     117] = 32'h0f40206f;
        ram_cell[     118] = 32'h00d00093;
        ram_cell[     119] = 32'h00b00113;
        ram_cell[     120] = 32'h002080b3;
        ram_cell[     121] = 32'h01800e93;
        ram_cell[     122] = 32'h01100193;
        ram_cell[     123] = 32'h01d08463;
        ram_cell[     124] = 32'h0d80206f;
        ram_cell[     125] = 32'h00e00093;
        ram_cell[     126] = 32'h00b00113;
        ram_cell[     127] = 32'h00208133;
        ram_cell[     128] = 32'h01900e93;
        ram_cell[     129] = 32'h01200193;
        ram_cell[     130] = 32'h01d10463;
        ram_cell[     131] = 32'h0bc0206f;
        ram_cell[     132] = 32'h00d00093;
        ram_cell[     133] = 32'h001080b3;
        ram_cell[     134] = 32'h01a00e93;
        ram_cell[     135] = 32'h01300193;
        ram_cell[     136] = 32'h01d08463;
        ram_cell[     137] = 32'h0a40206f;
        ram_cell[     138] = 32'h00000213;
        ram_cell[     139] = 32'h00d00093;
        ram_cell[     140] = 32'h00b00113;
        ram_cell[     141] = 32'h00208f33;
        ram_cell[     142] = 32'h000f0313;
        ram_cell[     143] = 32'h00120213;
        ram_cell[     144] = 32'h00200293;
        ram_cell[     145] = 32'hfe5214e3;
        ram_cell[     146] = 32'h01800e93;
        ram_cell[     147] = 32'h01400193;
        ram_cell[     148] = 32'h01d30463;
        ram_cell[     149] = 32'h0740206f;
        ram_cell[     150] = 32'h00000213;
        ram_cell[     151] = 32'h00e00093;
        ram_cell[     152] = 32'h00b00113;
        ram_cell[     153] = 32'h00208f33;
        ram_cell[     154] = 32'h00000013;
        ram_cell[     155] = 32'h000f0313;
        ram_cell[     156] = 32'h00120213;
        ram_cell[     157] = 32'h00200293;
        ram_cell[     158] = 32'hfe5212e3;
        ram_cell[     159] = 32'h01900e93;
        ram_cell[     160] = 32'h01500193;
        ram_cell[     161] = 32'h01d30463;
        ram_cell[     162] = 32'h0400206f;
        ram_cell[     163] = 32'h00000213;
        ram_cell[     164] = 32'h00f00093;
        ram_cell[     165] = 32'h00b00113;
        ram_cell[     166] = 32'h00208f33;
        ram_cell[     167] = 32'h00000013;
        ram_cell[     168] = 32'h00000013;
        ram_cell[     169] = 32'h000f0313;
        ram_cell[     170] = 32'h00120213;
        ram_cell[     171] = 32'h00200293;
        ram_cell[     172] = 32'hfe5210e3;
        ram_cell[     173] = 32'h01a00e93;
        ram_cell[     174] = 32'h01600193;
        ram_cell[     175] = 32'h01d30463;
        ram_cell[     176] = 32'h0080206f;
        ram_cell[     177] = 32'h00000213;
        ram_cell[     178] = 32'h00d00093;
        ram_cell[     179] = 32'h00b00113;
        ram_cell[     180] = 32'h00208f33;
        ram_cell[     181] = 32'h00120213;
        ram_cell[     182] = 32'h00200293;
        ram_cell[     183] = 32'hfe5216e3;
        ram_cell[     184] = 32'h01800e93;
        ram_cell[     185] = 32'h01700193;
        ram_cell[     186] = 32'h01df0463;
        ram_cell[     187] = 32'h7dd0106f;
        ram_cell[     188] = 32'h00000213;
        ram_cell[     189] = 32'h00e00093;
        ram_cell[     190] = 32'h00b00113;
        ram_cell[     191] = 32'h00000013;
        ram_cell[     192] = 32'h00208f33;
        ram_cell[     193] = 32'h00120213;
        ram_cell[     194] = 32'h00200293;
        ram_cell[     195] = 32'hfe5214e3;
        ram_cell[     196] = 32'h01900e93;
        ram_cell[     197] = 32'h01800193;
        ram_cell[     198] = 32'h01df0463;
        ram_cell[     199] = 32'h7ad0106f;
        ram_cell[     200] = 32'h00000213;
        ram_cell[     201] = 32'h00f00093;
        ram_cell[     202] = 32'h00b00113;
        ram_cell[     203] = 32'h00000013;
        ram_cell[     204] = 32'h00000013;
        ram_cell[     205] = 32'h00208f33;
        ram_cell[     206] = 32'h00120213;
        ram_cell[     207] = 32'h00200293;
        ram_cell[     208] = 32'hfe5212e3;
        ram_cell[     209] = 32'h01a00e93;
        ram_cell[     210] = 32'h01900193;
        ram_cell[     211] = 32'h01df0463;
        ram_cell[     212] = 32'h7790106f;
        ram_cell[     213] = 32'h00000213;
        ram_cell[     214] = 32'h00d00093;
        ram_cell[     215] = 32'h00000013;
        ram_cell[     216] = 32'h00b00113;
        ram_cell[     217] = 32'h00208f33;
        ram_cell[     218] = 32'h00120213;
        ram_cell[     219] = 32'h00200293;
        ram_cell[     220] = 32'hfe5214e3;
        ram_cell[     221] = 32'h01800e93;
        ram_cell[     222] = 32'h01a00193;
        ram_cell[     223] = 32'h01df0463;
        ram_cell[     224] = 32'h7490106f;
        ram_cell[     225] = 32'h00000213;
        ram_cell[     226] = 32'h00e00093;
        ram_cell[     227] = 32'h00000013;
        ram_cell[     228] = 32'h00b00113;
        ram_cell[     229] = 32'h00000013;
        ram_cell[     230] = 32'h00208f33;
        ram_cell[     231] = 32'h00120213;
        ram_cell[     232] = 32'h00200293;
        ram_cell[     233] = 32'hfe5212e3;
        ram_cell[     234] = 32'h01900e93;
        ram_cell[     235] = 32'h01b00193;
        ram_cell[     236] = 32'h01df0463;
        ram_cell[     237] = 32'h7150106f;
        ram_cell[     238] = 32'h00000213;
        ram_cell[     239] = 32'h00f00093;
        ram_cell[     240] = 32'h00000013;
        ram_cell[     241] = 32'h00000013;
        ram_cell[     242] = 32'h00b00113;
        ram_cell[     243] = 32'h00208f33;
        ram_cell[     244] = 32'h00120213;
        ram_cell[     245] = 32'h00200293;
        ram_cell[     246] = 32'hfe5212e3;
        ram_cell[     247] = 32'h01a00e93;
        ram_cell[     248] = 32'h01c00193;
        ram_cell[     249] = 32'h01df0463;
        ram_cell[     250] = 32'h6e10106f;
        ram_cell[     251] = 32'h00000213;
        ram_cell[     252] = 32'h00b00113;
        ram_cell[     253] = 32'h00d00093;
        ram_cell[     254] = 32'h00208f33;
        ram_cell[     255] = 32'h00120213;
        ram_cell[     256] = 32'h00200293;
        ram_cell[     257] = 32'hfe5216e3;
        ram_cell[     258] = 32'h01800e93;
        ram_cell[     259] = 32'h01d00193;
        ram_cell[     260] = 32'h01df0463;
        ram_cell[     261] = 32'h6b50106f;
        ram_cell[     262] = 32'h00000213;
        ram_cell[     263] = 32'h00b00113;
        ram_cell[     264] = 32'h00e00093;
        ram_cell[     265] = 32'h00000013;
        ram_cell[     266] = 32'h00208f33;
        ram_cell[     267] = 32'h00120213;
        ram_cell[     268] = 32'h00200293;
        ram_cell[     269] = 32'hfe5214e3;
        ram_cell[     270] = 32'h01900e93;
        ram_cell[     271] = 32'h01e00193;
        ram_cell[     272] = 32'h01df0463;
        ram_cell[     273] = 32'h6850106f;
        ram_cell[     274] = 32'h00000213;
        ram_cell[     275] = 32'h00b00113;
        ram_cell[     276] = 32'h00f00093;
        ram_cell[     277] = 32'h00000013;
        ram_cell[     278] = 32'h00000013;
        ram_cell[     279] = 32'h00208f33;
        ram_cell[     280] = 32'h00120213;
        ram_cell[     281] = 32'h00200293;
        ram_cell[     282] = 32'hfe5212e3;
        ram_cell[     283] = 32'h01a00e93;
        ram_cell[     284] = 32'h01f00193;
        ram_cell[     285] = 32'h01df0463;
        ram_cell[     286] = 32'h6510106f;
        ram_cell[     287] = 32'h00000213;
        ram_cell[     288] = 32'h00b00113;
        ram_cell[     289] = 32'h00000013;
        ram_cell[     290] = 32'h00d00093;
        ram_cell[     291] = 32'h00208f33;
        ram_cell[     292] = 32'h00120213;
        ram_cell[     293] = 32'h00200293;
        ram_cell[     294] = 32'hfe5214e3;
        ram_cell[     295] = 32'h01800e93;
        ram_cell[     296] = 32'h02000193;
        ram_cell[     297] = 32'h01df0463;
        ram_cell[     298] = 32'h6210106f;
        ram_cell[     299] = 32'h00000213;
        ram_cell[     300] = 32'h00b00113;
        ram_cell[     301] = 32'h00000013;
        ram_cell[     302] = 32'h00e00093;
        ram_cell[     303] = 32'h00000013;
        ram_cell[     304] = 32'h00208f33;
        ram_cell[     305] = 32'h00120213;
        ram_cell[     306] = 32'h00200293;
        ram_cell[     307] = 32'hfe5212e3;
        ram_cell[     308] = 32'h01900e93;
        ram_cell[     309] = 32'h02100193;
        ram_cell[     310] = 32'h01df0463;
        ram_cell[     311] = 32'h5ed0106f;
        ram_cell[     312] = 32'h00000213;
        ram_cell[     313] = 32'h00b00113;
        ram_cell[     314] = 32'h00000013;
        ram_cell[     315] = 32'h00000013;
        ram_cell[     316] = 32'h00f00093;
        ram_cell[     317] = 32'h00208f33;
        ram_cell[     318] = 32'h00120213;
        ram_cell[     319] = 32'h00200293;
        ram_cell[     320] = 32'hfe5212e3;
        ram_cell[     321] = 32'h01a00e93;
        ram_cell[     322] = 32'h02200193;
        ram_cell[     323] = 32'h01df0463;
        ram_cell[     324] = 32'h5b90106f;
        ram_cell[     325] = 32'h00f00093;
        ram_cell[     326] = 32'h00100133;
        ram_cell[     327] = 32'h00f00e93;
        ram_cell[     328] = 32'h02300193;
        ram_cell[     329] = 32'h01d10463;
        ram_cell[     330] = 32'h5a10106f;
        ram_cell[     331] = 32'h02000093;
        ram_cell[     332] = 32'h00008133;
        ram_cell[     333] = 32'h02000e93;
        ram_cell[     334] = 32'h02400193;
        ram_cell[     335] = 32'h01d10463;
        ram_cell[     336] = 32'h5890106f;
        ram_cell[     337] = 32'h000000b3;
        ram_cell[     338] = 32'h00000e93;
        ram_cell[     339] = 32'h02500193;
        ram_cell[     340] = 32'h01d08463;
        ram_cell[     341] = 32'h5750106f;
        ram_cell[     342] = 32'h01000093;
        ram_cell[     343] = 32'h01e00113;
        ram_cell[     344] = 32'h00208033;
        ram_cell[     345] = 32'h00000e93;
        ram_cell[     346] = 32'h02600193;
        ram_cell[     347] = 32'h01d00463;
        ram_cell[     348] = 32'h5590106f;
        ram_cell[     349] = 32'h00000093;
        ram_cell[     350] = 32'h00008f13;
        ram_cell[     351] = 32'h00000e93;
        ram_cell[     352] = 32'h02700193;
        ram_cell[     353] = 32'h01df0463;
        ram_cell[     354] = 32'h5410106f;
        ram_cell[     355] = 32'h00100093;
        ram_cell[     356] = 32'h00108f13;
        ram_cell[     357] = 32'h00200e93;
        ram_cell[     358] = 32'h02800193;
        ram_cell[     359] = 32'h01df0463;
        ram_cell[     360] = 32'h5290106f;
        ram_cell[     361] = 32'h00300093;
        ram_cell[     362] = 32'h00708f13;
        ram_cell[     363] = 32'h00a00e93;
        ram_cell[     364] = 32'h02900193;
        ram_cell[     365] = 32'h01df0463;
        ram_cell[     366] = 32'h5110106f;
        ram_cell[     367] = 32'h00000093;
        ram_cell[     368] = 32'h80008f13;
        ram_cell[     369] = 32'h80000e93;
        ram_cell[     370] = 32'h02a00193;
        ram_cell[     371] = 32'h01df0463;
        ram_cell[     372] = 32'h4f90106f;
        ram_cell[     373] = 32'h800000b7;
        ram_cell[     374] = 32'h00008f13;
        ram_cell[     375] = 32'h80000eb7;
        ram_cell[     376] = 32'h02b00193;
        ram_cell[     377] = 32'h01df0463;
        ram_cell[     378] = 32'h4e10106f;
        ram_cell[     379] = 32'h800000b7;
        ram_cell[     380] = 32'h80008f13;
        ram_cell[     381] = 32'h80000eb7;
        ram_cell[     382] = 32'h800e8e93;
        ram_cell[     383] = 32'h02c00193;
        ram_cell[     384] = 32'h01df0463;
        ram_cell[     385] = 32'h4c50106f;
        ram_cell[     386] = 32'h00000093;
        ram_cell[     387] = 32'h7ff08f13;
        ram_cell[     388] = 32'h7ff00e93;
        ram_cell[     389] = 32'h02d00193;
        ram_cell[     390] = 32'h01df0463;
        ram_cell[     391] = 32'h4ad0106f;
        ram_cell[     392] = 32'h800000b7;
        ram_cell[     393] = 32'hfff08093;
        ram_cell[     394] = 32'h00008f13;
        ram_cell[     395] = 32'h80000eb7;
        ram_cell[     396] = 32'hfffe8e93;
        ram_cell[     397] = 32'h02e00193;
        ram_cell[     398] = 32'h01df0463;
        ram_cell[     399] = 32'h48d0106f;
        ram_cell[     400] = 32'h800000b7;
        ram_cell[     401] = 32'hfff08093;
        ram_cell[     402] = 32'h7ff08f13;
        ram_cell[     403] = 32'h80000eb7;
        ram_cell[     404] = 32'h7fee8e93;
        ram_cell[     405] = 32'h02f00193;
        ram_cell[     406] = 32'h01df0463;
        ram_cell[     407] = 32'h46d0106f;
        ram_cell[     408] = 32'h800000b7;
        ram_cell[     409] = 32'h7ff08f13;
        ram_cell[     410] = 32'h80000eb7;
        ram_cell[     411] = 32'h7ffe8e93;
        ram_cell[     412] = 32'h03000193;
        ram_cell[     413] = 32'h01df0463;
        ram_cell[     414] = 32'h4510106f;
        ram_cell[     415] = 32'h800000b7;
        ram_cell[     416] = 32'hfff08093;
        ram_cell[     417] = 32'h80008f13;
        ram_cell[     418] = 32'h7ffffeb7;
        ram_cell[     419] = 32'h7ffe8e93;
        ram_cell[     420] = 32'h03100193;
        ram_cell[     421] = 32'h01df0463;
        ram_cell[     422] = 32'h4310106f;
        ram_cell[     423] = 32'h00000093;
        ram_cell[     424] = 32'hfff08f13;
        ram_cell[     425] = 32'hfff00e93;
        ram_cell[     426] = 32'h03200193;
        ram_cell[     427] = 32'h01df0463;
        ram_cell[     428] = 32'h4190106f;
        ram_cell[     429] = 32'hfff00093;
        ram_cell[     430] = 32'h00108f13;
        ram_cell[     431] = 32'h00000e93;
        ram_cell[     432] = 32'h03300193;
        ram_cell[     433] = 32'h01df0463;
        ram_cell[     434] = 32'h4010106f;
        ram_cell[     435] = 32'hfff00093;
        ram_cell[     436] = 32'hfff08f13;
        ram_cell[     437] = 32'hffe00e93;
        ram_cell[     438] = 32'h03400193;
        ram_cell[     439] = 32'h01df0463;
        ram_cell[     440] = 32'h3e90106f;
        ram_cell[     441] = 32'h800000b7;
        ram_cell[     442] = 32'hfff08093;
        ram_cell[     443] = 32'h00108f13;
        ram_cell[     444] = 32'h80000eb7;
        ram_cell[     445] = 32'h03500193;
        ram_cell[     446] = 32'h01df0463;
        ram_cell[     447] = 32'h3cd0106f;
        ram_cell[     448] = 32'h00d00093;
        ram_cell[     449] = 32'h00b08093;
        ram_cell[     450] = 32'h01800e93;
        ram_cell[     451] = 32'h03600193;
        ram_cell[     452] = 32'h01d08463;
        ram_cell[     453] = 32'h3b50106f;
        ram_cell[     454] = 32'h00000213;
        ram_cell[     455] = 32'h00d00093;
        ram_cell[     456] = 32'h00b08f13;
        ram_cell[     457] = 32'h000f0313;
        ram_cell[     458] = 32'h00120213;
        ram_cell[     459] = 32'h00200293;
        ram_cell[     460] = 32'hfe5216e3;
        ram_cell[     461] = 32'h01800e93;
        ram_cell[     462] = 32'h03700193;
        ram_cell[     463] = 32'h01d30463;
        ram_cell[     464] = 32'h3890106f;
        ram_cell[     465] = 32'h00000213;
        ram_cell[     466] = 32'h00d00093;
        ram_cell[     467] = 32'h00a08f13;
        ram_cell[     468] = 32'h00000013;
        ram_cell[     469] = 32'h000f0313;
        ram_cell[     470] = 32'h00120213;
        ram_cell[     471] = 32'h00200293;
        ram_cell[     472] = 32'hfe5214e3;
        ram_cell[     473] = 32'h01700e93;
        ram_cell[     474] = 32'h03800193;
        ram_cell[     475] = 32'h01d30463;
        ram_cell[     476] = 32'h3590106f;
        ram_cell[     477] = 32'h00000213;
        ram_cell[     478] = 32'h00d00093;
        ram_cell[     479] = 32'h00908f13;
        ram_cell[     480] = 32'h00000013;
        ram_cell[     481] = 32'h00000013;
        ram_cell[     482] = 32'h000f0313;
        ram_cell[     483] = 32'h00120213;
        ram_cell[     484] = 32'h00200293;
        ram_cell[     485] = 32'hfe5212e3;
        ram_cell[     486] = 32'h01600e93;
        ram_cell[     487] = 32'h03900193;
        ram_cell[     488] = 32'h01d30463;
        ram_cell[     489] = 32'h3250106f;
        ram_cell[     490] = 32'h00000213;
        ram_cell[     491] = 32'h00d00093;
        ram_cell[     492] = 32'h00b08f13;
        ram_cell[     493] = 32'h00120213;
        ram_cell[     494] = 32'h00200293;
        ram_cell[     495] = 32'hfe5218e3;
        ram_cell[     496] = 32'h01800e93;
        ram_cell[     497] = 32'h03a00193;
        ram_cell[     498] = 32'h01df0463;
        ram_cell[     499] = 32'h2fd0106f;
        ram_cell[     500] = 32'h00000213;
        ram_cell[     501] = 32'h00d00093;
        ram_cell[     502] = 32'h00000013;
        ram_cell[     503] = 32'h00a08f13;
        ram_cell[     504] = 32'h00120213;
        ram_cell[     505] = 32'h00200293;
        ram_cell[     506] = 32'hfe5216e3;
        ram_cell[     507] = 32'h01700e93;
        ram_cell[     508] = 32'h03b00193;
        ram_cell[     509] = 32'h01df0463;
        ram_cell[     510] = 32'h2d10106f;
        ram_cell[     511] = 32'h00000213;
        ram_cell[     512] = 32'h00d00093;
        ram_cell[     513] = 32'h00000013;
        ram_cell[     514] = 32'h00000013;
        ram_cell[     515] = 32'h00908f13;
        ram_cell[     516] = 32'h00120213;
        ram_cell[     517] = 32'h00200293;
        ram_cell[     518] = 32'hfe5214e3;
        ram_cell[     519] = 32'h01600e93;
        ram_cell[     520] = 32'h03c00193;
        ram_cell[     521] = 32'h01df0463;
        ram_cell[     522] = 32'h2a10106f;
        ram_cell[     523] = 32'h02000093;
        ram_cell[     524] = 32'h02000e93;
        ram_cell[     525] = 32'h03d00193;
        ram_cell[     526] = 32'h01d08463;
        ram_cell[     527] = 32'h28d0106f;
        ram_cell[     528] = 32'h02100093;
        ram_cell[     529] = 32'h03208013;
        ram_cell[     530] = 32'h00000e93;
        ram_cell[     531] = 32'h03e00193;
        ram_cell[     532] = 32'h01d00463;
        ram_cell[     533] = 32'h2750106f;
        ram_cell[     534] = 32'hff0100b7;
        ram_cell[     535] = 32'hf0008093;
        ram_cell[     536] = 32'h0f0f1137;
        ram_cell[     537] = 32'hf0f10113;
        ram_cell[     538] = 32'h0020ff33;
        ram_cell[     539] = 32'h0f001eb7;
        ram_cell[     540] = 32'hf00e8e93;
        ram_cell[     541] = 32'h03f00193;
        ram_cell[     542] = 32'h01df0463;
        ram_cell[     543] = 32'h24d0106f;
        ram_cell[     544] = 32'h0ff010b7;
        ram_cell[     545] = 32'hff008093;
        ram_cell[     546] = 32'hf0f0f137;
        ram_cell[     547] = 32'h0f010113;
        ram_cell[     548] = 32'h0020ff33;
        ram_cell[     549] = 32'h00f00eb7;
        ram_cell[     550] = 32'h0f0e8e93;
        ram_cell[     551] = 32'h04000193;
        ram_cell[     552] = 32'h01df0463;
        ram_cell[     553] = 32'h2250106f;
        ram_cell[     554] = 32'h00ff00b7;
        ram_cell[     555] = 32'h0ff08093;
        ram_cell[     556] = 32'h0f0f1137;
        ram_cell[     557] = 32'hf0f10113;
        ram_cell[     558] = 32'h0020ff33;
        ram_cell[     559] = 32'h000f0eb7;
        ram_cell[     560] = 32'h00fe8e93;
        ram_cell[     561] = 32'h04100193;
        ram_cell[     562] = 32'h01df0463;
        ram_cell[     563] = 32'h1fd0106f;
        ram_cell[     564] = 32'hf00ff0b7;
        ram_cell[     565] = 32'h00f08093;
        ram_cell[     566] = 32'hf0f0f137;
        ram_cell[     567] = 32'h0f010113;
        ram_cell[     568] = 32'h0020ff33;
        ram_cell[     569] = 32'hf000feb7;
        ram_cell[     570] = 32'h04200193;
        ram_cell[     571] = 32'h01df0463;
        ram_cell[     572] = 32'h1d90106f;
        ram_cell[     573] = 32'hff0100b7;
        ram_cell[     574] = 32'hf0008093;
        ram_cell[     575] = 32'h0f0f1137;
        ram_cell[     576] = 32'hf0f10113;
        ram_cell[     577] = 32'h0020f0b3;
        ram_cell[     578] = 32'h0f001eb7;
        ram_cell[     579] = 32'hf00e8e93;
        ram_cell[     580] = 32'h04300193;
        ram_cell[     581] = 32'h01d08463;
        ram_cell[     582] = 32'h1b10106f;
        ram_cell[     583] = 32'h0ff010b7;
        ram_cell[     584] = 32'hff008093;
        ram_cell[     585] = 32'hf0f0f137;
        ram_cell[     586] = 32'h0f010113;
        ram_cell[     587] = 32'h0020f133;
        ram_cell[     588] = 32'h00f00eb7;
        ram_cell[     589] = 32'h0f0e8e93;
        ram_cell[     590] = 32'h04400193;
        ram_cell[     591] = 32'h01d10463;
        ram_cell[     592] = 32'h1890106f;
        ram_cell[     593] = 32'hff0100b7;
        ram_cell[     594] = 32'hf0008093;
        ram_cell[     595] = 32'h0010f0b3;
        ram_cell[     596] = 32'hff010eb7;
        ram_cell[     597] = 32'hf00e8e93;
        ram_cell[     598] = 32'h04500193;
        ram_cell[     599] = 32'h01d08463;
        ram_cell[     600] = 32'h1690106f;
        ram_cell[     601] = 32'h00000213;
        ram_cell[     602] = 32'hff0100b7;
        ram_cell[     603] = 32'hf0008093;
        ram_cell[     604] = 32'h0f0f1137;
        ram_cell[     605] = 32'hf0f10113;
        ram_cell[     606] = 32'h0020ff33;
        ram_cell[     607] = 32'h000f0313;
        ram_cell[     608] = 32'h00120213;
        ram_cell[     609] = 32'h00200293;
        ram_cell[     610] = 32'hfe5210e3;
        ram_cell[     611] = 32'h0f001eb7;
        ram_cell[     612] = 32'hf00e8e93;
        ram_cell[     613] = 32'h04600193;
        ram_cell[     614] = 32'h01d30463;
        ram_cell[     615] = 32'h12d0106f;
        ram_cell[     616] = 32'h00000213;
        ram_cell[     617] = 32'h0ff010b7;
        ram_cell[     618] = 32'hff008093;
        ram_cell[     619] = 32'hf0f0f137;
        ram_cell[     620] = 32'h0f010113;
        ram_cell[     621] = 32'h0020ff33;
        ram_cell[     622] = 32'h00000013;
        ram_cell[     623] = 32'h000f0313;
        ram_cell[     624] = 32'h00120213;
        ram_cell[     625] = 32'h00200293;
        ram_cell[     626] = 32'hfc521ee3;
        ram_cell[     627] = 32'h00f00eb7;
        ram_cell[     628] = 32'h0f0e8e93;
        ram_cell[     629] = 32'h04700193;
        ram_cell[     630] = 32'h01d30463;
        ram_cell[     631] = 32'h0ed0106f;
        ram_cell[     632] = 32'h00000213;
        ram_cell[     633] = 32'h00ff00b7;
        ram_cell[     634] = 32'h0ff08093;
        ram_cell[     635] = 32'h0f0f1137;
        ram_cell[     636] = 32'hf0f10113;
        ram_cell[     637] = 32'h0020ff33;
        ram_cell[     638] = 32'h00000013;
        ram_cell[     639] = 32'h00000013;
        ram_cell[     640] = 32'h000f0313;
        ram_cell[     641] = 32'h00120213;
        ram_cell[     642] = 32'h00200293;
        ram_cell[     643] = 32'hfc521ce3;
        ram_cell[     644] = 32'h000f0eb7;
        ram_cell[     645] = 32'h00fe8e93;
        ram_cell[     646] = 32'h04800193;
        ram_cell[     647] = 32'h01d30463;
        ram_cell[     648] = 32'h0a90106f;
        ram_cell[     649] = 32'h00000213;
        ram_cell[     650] = 32'hff0100b7;
        ram_cell[     651] = 32'hf0008093;
        ram_cell[     652] = 32'h0f0f1137;
        ram_cell[     653] = 32'hf0f10113;
        ram_cell[     654] = 32'h0020ff33;
        ram_cell[     655] = 32'h00120213;
        ram_cell[     656] = 32'h00200293;
        ram_cell[     657] = 32'hfe5212e3;
        ram_cell[     658] = 32'h0f001eb7;
        ram_cell[     659] = 32'hf00e8e93;
        ram_cell[     660] = 32'h04900193;
        ram_cell[     661] = 32'h01df0463;
        ram_cell[     662] = 32'h0710106f;
        ram_cell[     663] = 32'h00000213;
        ram_cell[     664] = 32'h0ff010b7;
        ram_cell[     665] = 32'hff008093;
        ram_cell[     666] = 32'hf0f0f137;
        ram_cell[     667] = 32'h0f010113;
        ram_cell[     668] = 32'h00000013;
        ram_cell[     669] = 32'h0020ff33;
        ram_cell[     670] = 32'h00120213;
        ram_cell[     671] = 32'h00200293;
        ram_cell[     672] = 32'hfe5210e3;
        ram_cell[     673] = 32'h00f00eb7;
        ram_cell[     674] = 32'h0f0e8e93;
        ram_cell[     675] = 32'h04a00193;
        ram_cell[     676] = 32'h01df0463;
        ram_cell[     677] = 32'h0350106f;
        ram_cell[     678] = 32'h00000213;
        ram_cell[     679] = 32'h00ff00b7;
        ram_cell[     680] = 32'h0ff08093;
        ram_cell[     681] = 32'h0f0f1137;
        ram_cell[     682] = 32'hf0f10113;
        ram_cell[     683] = 32'h00000013;
        ram_cell[     684] = 32'h00000013;
        ram_cell[     685] = 32'h0020ff33;
        ram_cell[     686] = 32'h00120213;
        ram_cell[     687] = 32'h00200293;
        ram_cell[     688] = 32'hfc521ee3;
        ram_cell[     689] = 32'h000f0eb7;
        ram_cell[     690] = 32'h00fe8e93;
        ram_cell[     691] = 32'h04b00193;
        ram_cell[     692] = 32'h01df0463;
        ram_cell[     693] = 32'h7f40106f;
        ram_cell[     694] = 32'h00000213;
        ram_cell[     695] = 32'hff0100b7;
        ram_cell[     696] = 32'hf0008093;
        ram_cell[     697] = 32'h00000013;
        ram_cell[     698] = 32'h0f0f1137;
        ram_cell[     699] = 32'hf0f10113;
        ram_cell[     700] = 32'h0020ff33;
        ram_cell[     701] = 32'h00120213;
        ram_cell[     702] = 32'h00200293;
        ram_cell[     703] = 32'hfe5210e3;
        ram_cell[     704] = 32'h0f001eb7;
        ram_cell[     705] = 32'hf00e8e93;
        ram_cell[     706] = 32'h04c00193;
        ram_cell[     707] = 32'h01df0463;
        ram_cell[     708] = 32'h7b80106f;
        ram_cell[     709] = 32'h00000213;
        ram_cell[     710] = 32'h0ff010b7;
        ram_cell[     711] = 32'hff008093;
        ram_cell[     712] = 32'h00000013;
        ram_cell[     713] = 32'hf0f0f137;
        ram_cell[     714] = 32'h0f010113;
        ram_cell[     715] = 32'h00000013;
        ram_cell[     716] = 32'h0020ff33;
        ram_cell[     717] = 32'h00120213;
        ram_cell[     718] = 32'h00200293;
        ram_cell[     719] = 32'hfc521ee3;
        ram_cell[     720] = 32'h00f00eb7;
        ram_cell[     721] = 32'h0f0e8e93;
        ram_cell[     722] = 32'h04d00193;
        ram_cell[     723] = 32'h01df0463;
        ram_cell[     724] = 32'h7780106f;
        ram_cell[     725] = 32'h00000213;
        ram_cell[     726] = 32'h00ff00b7;
        ram_cell[     727] = 32'h0ff08093;
        ram_cell[     728] = 32'h00000013;
        ram_cell[     729] = 32'h00000013;
        ram_cell[     730] = 32'h0f0f1137;
        ram_cell[     731] = 32'hf0f10113;
        ram_cell[     732] = 32'h0020ff33;
        ram_cell[     733] = 32'h00120213;
        ram_cell[     734] = 32'h00200293;
        ram_cell[     735] = 32'hfc521ee3;
        ram_cell[     736] = 32'h000f0eb7;
        ram_cell[     737] = 32'h00fe8e93;
        ram_cell[     738] = 32'h04e00193;
        ram_cell[     739] = 32'h01df0463;
        ram_cell[     740] = 32'h7380106f;
        ram_cell[     741] = 32'h00000213;
        ram_cell[     742] = 32'h0f0f1137;
        ram_cell[     743] = 32'hf0f10113;
        ram_cell[     744] = 32'hff0100b7;
        ram_cell[     745] = 32'hf0008093;
        ram_cell[     746] = 32'h0020ff33;
        ram_cell[     747] = 32'h00120213;
        ram_cell[     748] = 32'h00200293;
        ram_cell[     749] = 32'hfe5212e3;
        ram_cell[     750] = 32'h0f001eb7;
        ram_cell[     751] = 32'hf00e8e93;
        ram_cell[     752] = 32'h04f00193;
        ram_cell[     753] = 32'h01df0463;
        ram_cell[     754] = 32'h7000106f;
        ram_cell[     755] = 32'h00000213;
        ram_cell[     756] = 32'hf0f0f137;
        ram_cell[     757] = 32'h0f010113;
        ram_cell[     758] = 32'h0ff010b7;
        ram_cell[     759] = 32'hff008093;
        ram_cell[     760] = 32'h00000013;
        ram_cell[     761] = 32'h0020ff33;
        ram_cell[     762] = 32'h00120213;
        ram_cell[     763] = 32'h00200293;
        ram_cell[     764] = 32'hfe5210e3;
        ram_cell[     765] = 32'h00f00eb7;
        ram_cell[     766] = 32'h0f0e8e93;
        ram_cell[     767] = 32'h05000193;
        ram_cell[     768] = 32'h01df0463;
        ram_cell[     769] = 32'h6c40106f;
        ram_cell[     770] = 32'h00000213;
        ram_cell[     771] = 32'h0f0f1137;
        ram_cell[     772] = 32'hf0f10113;
        ram_cell[     773] = 32'h00ff00b7;
        ram_cell[     774] = 32'h0ff08093;
        ram_cell[     775] = 32'h00000013;
        ram_cell[     776] = 32'h00000013;
        ram_cell[     777] = 32'h0020ff33;
        ram_cell[     778] = 32'h00120213;
        ram_cell[     779] = 32'h00200293;
        ram_cell[     780] = 32'hfc521ee3;
        ram_cell[     781] = 32'h000f0eb7;
        ram_cell[     782] = 32'h00fe8e93;
        ram_cell[     783] = 32'h05100193;
        ram_cell[     784] = 32'h01df0463;
        ram_cell[     785] = 32'h6840106f;
        ram_cell[     786] = 32'h00000213;
        ram_cell[     787] = 32'h0f0f1137;
        ram_cell[     788] = 32'hf0f10113;
        ram_cell[     789] = 32'h00000013;
        ram_cell[     790] = 32'hff0100b7;
        ram_cell[     791] = 32'hf0008093;
        ram_cell[     792] = 32'h0020ff33;
        ram_cell[     793] = 32'h00120213;
        ram_cell[     794] = 32'h00200293;
        ram_cell[     795] = 32'hfe5210e3;
        ram_cell[     796] = 32'h0f001eb7;
        ram_cell[     797] = 32'hf00e8e93;
        ram_cell[     798] = 32'h05200193;
        ram_cell[     799] = 32'h01df0463;
        ram_cell[     800] = 32'h6480106f;
        ram_cell[     801] = 32'h00000213;
        ram_cell[     802] = 32'hf0f0f137;
        ram_cell[     803] = 32'h0f010113;
        ram_cell[     804] = 32'h00000013;
        ram_cell[     805] = 32'h0ff010b7;
        ram_cell[     806] = 32'hff008093;
        ram_cell[     807] = 32'h00000013;
        ram_cell[     808] = 32'h0020ff33;
        ram_cell[     809] = 32'h00120213;
        ram_cell[     810] = 32'h00200293;
        ram_cell[     811] = 32'hfc521ee3;
        ram_cell[     812] = 32'h00f00eb7;
        ram_cell[     813] = 32'h0f0e8e93;
        ram_cell[     814] = 32'h05300193;
        ram_cell[     815] = 32'h01df0463;
        ram_cell[     816] = 32'h6080106f;
        ram_cell[     817] = 32'h00000213;
        ram_cell[     818] = 32'h0f0f1137;
        ram_cell[     819] = 32'hf0f10113;
        ram_cell[     820] = 32'h00000013;
        ram_cell[     821] = 32'h00000013;
        ram_cell[     822] = 32'h00ff00b7;
        ram_cell[     823] = 32'h0ff08093;
        ram_cell[     824] = 32'h0020ff33;
        ram_cell[     825] = 32'h00120213;
        ram_cell[     826] = 32'h00200293;
        ram_cell[     827] = 32'hfc521ee3;
        ram_cell[     828] = 32'h000f0eb7;
        ram_cell[     829] = 32'h00fe8e93;
        ram_cell[     830] = 32'h05400193;
        ram_cell[     831] = 32'h01df0463;
        ram_cell[     832] = 32'h5c80106f;
        ram_cell[     833] = 32'hff0100b7;
        ram_cell[     834] = 32'hf0008093;
        ram_cell[     835] = 32'h00107133;
        ram_cell[     836] = 32'h00000e93;
        ram_cell[     837] = 32'h05500193;
        ram_cell[     838] = 32'h01d10463;
        ram_cell[     839] = 32'h5ac0106f;
        ram_cell[     840] = 32'h00ff00b7;
        ram_cell[     841] = 32'h0ff08093;
        ram_cell[     842] = 32'h0000f133;
        ram_cell[     843] = 32'h00000e93;
        ram_cell[     844] = 32'h05600193;
        ram_cell[     845] = 32'h01d10463;
        ram_cell[     846] = 32'h5900106f;
        ram_cell[     847] = 32'h000070b3;
        ram_cell[     848] = 32'h00000e93;
        ram_cell[     849] = 32'h05700193;
        ram_cell[     850] = 32'h01d08463;
        ram_cell[     851] = 32'h57c0106f;
        ram_cell[     852] = 32'h111110b7;
        ram_cell[     853] = 32'h11108093;
        ram_cell[     854] = 32'h22222137;
        ram_cell[     855] = 32'h22210113;
        ram_cell[     856] = 32'h0020f033;
        ram_cell[     857] = 32'h00000e93;
        ram_cell[     858] = 32'h05800193;
        ram_cell[     859] = 32'h01d00463;
        ram_cell[     860] = 32'h5580106f;
        ram_cell[     861] = 32'hff0100b7;
        ram_cell[     862] = 32'hf0008093;
        ram_cell[     863] = 32'hf0f0ff13;
        ram_cell[     864] = 32'hff010eb7;
        ram_cell[     865] = 32'hf00e8e93;
        ram_cell[     866] = 32'h05900193;
        ram_cell[     867] = 32'h01df0463;
        ram_cell[     868] = 32'h5380106f;
        ram_cell[     869] = 32'h0ff010b7;
        ram_cell[     870] = 32'hff008093;
        ram_cell[     871] = 32'h0f00ff13;
        ram_cell[     872] = 32'h0f000e93;
        ram_cell[     873] = 32'h05a00193;
        ram_cell[     874] = 32'h01df0463;
        ram_cell[     875] = 32'h51c0106f;
        ram_cell[     876] = 32'h00ff00b7;
        ram_cell[     877] = 32'h0ff08093;
        ram_cell[     878] = 32'h70f0ff13;
        ram_cell[     879] = 32'h00f00e93;
        ram_cell[     880] = 32'h05b00193;
        ram_cell[     881] = 32'h01df0463;
        ram_cell[     882] = 32'h5000106f;
        ram_cell[     883] = 32'hf00ff0b7;
        ram_cell[     884] = 32'h00f08093;
        ram_cell[     885] = 32'h0f00ff13;
        ram_cell[     886] = 32'h00000e93;
        ram_cell[     887] = 32'h05c00193;
        ram_cell[     888] = 32'h01df0463;
        ram_cell[     889] = 32'h4e40106f;
        ram_cell[     890] = 32'hff0100b7;
        ram_cell[     891] = 32'hf0008093;
        ram_cell[     892] = 32'h0f00f093;
        ram_cell[     893] = 32'h00000e93;
        ram_cell[     894] = 32'h05d00193;
        ram_cell[     895] = 32'h01d08463;
        ram_cell[     896] = 32'h4c80106f;
        ram_cell[     897] = 32'h00000213;
        ram_cell[     898] = 32'h0ff010b7;
        ram_cell[     899] = 32'hff008093;
        ram_cell[     900] = 32'h70f0ff13;
        ram_cell[     901] = 32'h000f0313;
        ram_cell[     902] = 32'h00120213;
        ram_cell[     903] = 32'h00200293;
        ram_cell[     904] = 32'hfe5214e3;
        ram_cell[     905] = 32'h70000e93;
        ram_cell[     906] = 32'h05e00193;
        ram_cell[     907] = 32'h01d30463;
        ram_cell[     908] = 32'h4980106f;
        ram_cell[     909] = 32'h00000213;
        ram_cell[     910] = 32'h00ff00b7;
        ram_cell[     911] = 32'h0ff08093;
        ram_cell[     912] = 32'h0f00ff13;
        ram_cell[     913] = 32'h00000013;
        ram_cell[     914] = 32'h000f0313;
        ram_cell[     915] = 32'h00120213;
        ram_cell[     916] = 32'h00200293;
        ram_cell[     917] = 32'hfe5212e3;
        ram_cell[     918] = 32'h0f000e93;
        ram_cell[     919] = 32'h05f00193;
        ram_cell[     920] = 32'h01d30463;
        ram_cell[     921] = 32'h4640106f;
        ram_cell[     922] = 32'h00000213;
        ram_cell[     923] = 32'hf00ff0b7;
        ram_cell[     924] = 32'h00f08093;
        ram_cell[     925] = 32'hf0f0ff13;
        ram_cell[     926] = 32'h00000013;
        ram_cell[     927] = 32'h00000013;
        ram_cell[     928] = 32'h000f0313;
        ram_cell[     929] = 32'h00120213;
        ram_cell[     930] = 32'h00200293;
        ram_cell[     931] = 32'hfe5210e3;
        ram_cell[     932] = 32'hf00ffeb7;
        ram_cell[     933] = 32'h00fe8e93;
        ram_cell[     934] = 32'h06000193;
        ram_cell[     935] = 32'h01d30463;
        ram_cell[     936] = 32'h4280106f;
        ram_cell[     937] = 32'h00000213;
        ram_cell[     938] = 32'h0ff010b7;
        ram_cell[     939] = 32'hff008093;
        ram_cell[     940] = 32'h70f0ff13;
        ram_cell[     941] = 32'h00120213;
        ram_cell[     942] = 32'h00200293;
        ram_cell[     943] = 32'hfe5216e3;
        ram_cell[     944] = 32'h70000e93;
        ram_cell[     945] = 32'h06100193;
        ram_cell[     946] = 32'h01df0463;
        ram_cell[     947] = 32'h3fc0106f;
        ram_cell[     948] = 32'h00000213;
        ram_cell[     949] = 32'h00ff00b7;
        ram_cell[     950] = 32'h0ff08093;
        ram_cell[     951] = 32'h00000013;
        ram_cell[     952] = 32'h0f00ff13;
        ram_cell[     953] = 32'h00120213;
        ram_cell[     954] = 32'h00200293;
        ram_cell[     955] = 32'hfe5214e3;
        ram_cell[     956] = 32'h0f000e93;
        ram_cell[     957] = 32'h06200193;
        ram_cell[     958] = 32'h01df0463;
        ram_cell[     959] = 32'h3cc0106f;
        ram_cell[     960] = 32'h00000213;
        ram_cell[     961] = 32'hf00ff0b7;
        ram_cell[     962] = 32'h00f08093;
        ram_cell[     963] = 32'h00000013;
        ram_cell[     964] = 32'h00000013;
        ram_cell[     965] = 32'h70f0ff13;
        ram_cell[     966] = 32'h00120213;
        ram_cell[     967] = 32'h00200293;
        ram_cell[     968] = 32'hfe5212e3;
        ram_cell[     969] = 32'h00f00e93;
        ram_cell[     970] = 32'h06300193;
        ram_cell[     971] = 32'h01df0463;
        ram_cell[     972] = 32'h3980106f;
        ram_cell[     973] = 32'h0f007093;
        ram_cell[     974] = 32'h00000e93;
        ram_cell[     975] = 32'h06400193;
        ram_cell[     976] = 32'h01d08463;
        ram_cell[     977] = 32'h3840106f;
        ram_cell[     978] = 32'h00ff00b7;
        ram_cell[     979] = 32'h0ff08093;
        ram_cell[     980] = 32'h70f0f013;
        ram_cell[     981] = 32'h00000e93;
        ram_cell[     982] = 32'h06500193;
        ram_cell[     983] = 32'h01d00463;
        ram_cell[     984] = 32'h3680106f;
        ram_cell[     985] = 32'h00000013;
        ram_cell[     986] = 32'h00002517;
        ram_cell[     987] = 32'h71c50513;
        ram_cell[     988] = 32'h004005ef;
        ram_cell[     989] = 32'h40b50533;
        ram_cell[     990] = 32'h00002eb7;
        ram_cell[     991] = 32'h710e8e93;
        ram_cell[     992] = 32'h06600193;
        ram_cell[     993] = 32'h01d50463;
        ram_cell[     994] = 32'h3400106f;
        ram_cell[     995] = 32'h00000013;
        ram_cell[     996] = 32'hffffe517;
        ram_cell[     997] = 32'h8fc50513;
        ram_cell[     998] = 32'h004005ef;
        ram_cell[     999] = 32'h40b50533;
        ram_cell[    1000] = 32'hffffeeb7;
        ram_cell[    1001] = 32'h8f0e8e93;
        ram_cell[    1002] = 32'h06700193;
        ram_cell[    1003] = 32'h01d50463;
        ram_cell[    1004] = 32'h3180106f;
        ram_cell[    1005] = 32'h06800193;
        ram_cell[    1006] = 32'h00000093;
        ram_cell[    1007] = 32'h00000113;
        ram_cell[    1008] = 32'h00208863;
        ram_cell[    1009] = 32'h00300463;
        ram_cell[    1010] = 32'h3000106f;
        ram_cell[    1011] = 32'h00301863;
        ram_cell[    1012] = 32'hfe208ee3;
        ram_cell[    1013] = 32'h00300463;
        ram_cell[    1014] = 32'h2f00106f;
        ram_cell[    1015] = 32'h06900193;
        ram_cell[    1016] = 32'h00100093;
        ram_cell[    1017] = 32'h00100113;
        ram_cell[    1018] = 32'h00208863;
        ram_cell[    1019] = 32'h00300463;
        ram_cell[    1020] = 32'h2d80106f;
        ram_cell[    1021] = 32'h00301863;
        ram_cell[    1022] = 32'hfe208ee3;
        ram_cell[    1023] = 32'h00300463;
        ram_cell[    1024] = 32'h2c80106f;
        ram_cell[    1025] = 32'h06a00193;
        ram_cell[    1026] = 32'hfff00093;
        ram_cell[    1027] = 32'hfff00113;
        ram_cell[    1028] = 32'h00208863;
        ram_cell[    1029] = 32'h00300463;
        ram_cell[    1030] = 32'h2b00106f;
        ram_cell[    1031] = 32'h00301863;
        ram_cell[    1032] = 32'hfe208ee3;
        ram_cell[    1033] = 32'h00300463;
        ram_cell[    1034] = 32'h2a00106f;
        ram_cell[    1035] = 32'h06b00193;
        ram_cell[    1036] = 32'h00000093;
        ram_cell[    1037] = 32'h00100113;
        ram_cell[    1038] = 32'h00208463;
        ram_cell[    1039] = 32'h00301663;
        ram_cell[    1040] = 32'h00300463;
        ram_cell[    1041] = 32'h2840106f;
        ram_cell[    1042] = 32'hfe208ce3;
        ram_cell[    1043] = 32'h06c00193;
        ram_cell[    1044] = 32'h00100093;
        ram_cell[    1045] = 32'h00000113;
        ram_cell[    1046] = 32'h00208463;
        ram_cell[    1047] = 32'h00301663;
        ram_cell[    1048] = 32'h00300463;
        ram_cell[    1049] = 32'h2640106f;
        ram_cell[    1050] = 32'hfe208ce3;
        ram_cell[    1051] = 32'h06d00193;
        ram_cell[    1052] = 32'hfff00093;
        ram_cell[    1053] = 32'h00100113;
        ram_cell[    1054] = 32'h00208463;
        ram_cell[    1055] = 32'h00301663;
        ram_cell[    1056] = 32'h00300463;
        ram_cell[    1057] = 32'h2440106f;
        ram_cell[    1058] = 32'hfe208ce3;
        ram_cell[    1059] = 32'h06e00193;
        ram_cell[    1060] = 32'h00100093;
        ram_cell[    1061] = 32'hfff00113;
        ram_cell[    1062] = 32'h00208463;
        ram_cell[    1063] = 32'h00301663;
        ram_cell[    1064] = 32'h00300463;
        ram_cell[    1065] = 32'h2240106f;
        ram_cell[    1066] = 32'hfe208ce3;
        ram_cell[    1067] = 32'h06f00193;
        ram_cell[    1068] = 32'h00000213;
        ram_cell[    1069] = 32'h00000093;
        ram_cell[    1070] = 32'hfff00113;
        ram_cell[    1071] = 32'h00209463;
        ram_cell[    1072] = 32'h2080106f;
        ram_cell[    1073] = 32'h00120213;
        ram_cell[    1074] = 32'h00200293;
        ram_cell[    1075] = 32'hfe5214e3;
        ram_cell[    1076] = 32'h07000193;
        ram_cell[    1077] = 32'h00000213;
        ram_cell[    1078] = 32'h00000093;
        ram_cell[    1079] = 32'hfff00113;
        ram_cell[    1080] = 32'h00000013;
        ram_cell[    1081] = 32'h00209463;
        ram_cell[    1082] = 32'h1e00106f;
        ram_cell[    1083] = 32'h00120213;
        ram_cell[    1084] = 32'h00200293;
        ram_cell[    1085] = 32'hfe5212e3;
        ram_cell[    1086] = 32'h07100193;
        ram_cell[    1087] = 32'h00000213;
        ram_cell[    1088] = 32'h00000093;
        ram_cell[    1089] = 32'hfff00113;
        ram_cell[    1090] = 32'h00000013;
        ram_cell[    1091] = 32'h00000013;
        ram_cell[    1092] = 32'h00209463;
        ram_cell[    1093] = 32'h1b40106f;
        ram_cell[    1094] = 32'h00120213;
        ram_cell[    1095] = 32'h00200293;
        ram_cell[    1096] = 32'hfe5210e3;
        ram_cell[    1097] = 32'h07200193;
        ram_cell[    1098] = 32'h00000213;
        ram_cell[    1099] = 32'h00000093;
        ram_cell[    1100] = 32'h00000013;
        ram_cell[    1101] = 32'hfff00113;
        ram_cell[    1102] = 32'h00209463;
        ram_cell[    1103] = 32'h18c0106f;
        ram_cell[    1104] = 32'h00120213;
        ram_cell[    1105] = 32'h00200293;
        ram_cell[    1106] = 32'hfe5212e3;
        ram_cell[    1107] = 32'h07300193;
        ram_cell[    1108] = 32'h00000213;
        ram_cell[    1109] = 32'h00000093;
        ram_cell[    1110] = 32'h00000013;
        ram_cell[    1111] = 32'hfff00113;
        ram_cell[    1112] = 32'h00000013;
        ram_cell[    1113] = 32'h00209463;
        ram_cell[    1114] = 32'h1600106f;
        ram_cell[    1115] = 32'h00120213;
        ram_cell[    1116] = 32'h00200293;
        ram_cell[    1117] = 32'hfe5210e3;
        ram_cell[    1118] = 32'h07400193;
        ram_cell[    1119] = 32'h00000213;
        ram_cell[    1120] = 32'h00000093;
        ram_cell[    1121] = 32'h00000013;
        ram_cell[    1122] = 32'h00000013;
        ram_cell[    1123] = 32'hfff00113;
        ram_cell[    1124] = 32'h00209463;
        ram_cell[    1125] = 32'h1340106f;
        ram_cell[    1126] = 32'h00120213;
        ram_cell[    1127] = 32'h00200293;
        ram_cell[    1128] = 32'hfe5210e3;
        ram_cell[    1129] = 32'h07500193;
        ram_cell[    1130] = 32'h00000213;
        ram_cell[    1131] = 32'h00000093;
        ram_cell[    1132] = 32'hfff00113;
        ram_cell[    1133] = 32'h00209463;
        ram_cell[    1134] = 32'h1100106f;
        ram_cell[    1135] = 32'h00120213;
        ram_cell[    1136] = 32'h00200293;
        ram_cell[    1137] = 32'hfe5214e3;
        ram_cell[    1138] = 32'h07600193;
        ram_cell[    1139] = 32'h00000213;
        ram_cell[    1140] = 32'h00000093;
        ram_cell[    1141] = 32'hfff00113;
        ram_cell[    1142] = 32'h00000013;
        ram_cell[    1143] = 32'h00209463;
        ram_cell[    1144] = 32'h0e80106f;
        ram_cell[    1145] = 32'h00120213;
        ram_cell[    1146] = 32'h00200293;
        ram_cell[    1147] = 32'hfe5212e3;
        ram_cell[    1148] = 32'h07700193;
        ram_cell[    1149] = 32'h00000213;
        ram_cell[    1150] = 32'h00000093;
        ram_cell[    1151] = 32'hfff00113;
        ram_cell[    1152] = 32'h00000013;
        ram_cell[    1153] = 32'h00000013;
        ram_cell[    1154] = 32'h00209463;
        ram_cell[    1155] = 32'h0bc0106f;
        ram_cell[    1156] = 32'h00120213;
        ram_cell[    1157] = 32'h00200293;
        ram_cell[    1158] = 32'hfe5210e3;
        ram_cell[    1159] = 32'h07800193;
        ram_cell[    1160] = 32'h00000213;
        ram_cell[    1161] = 32'h00000093;
        ram_cell[    1162] = 32'h00000013;
        ram_cell[    1163] = 32'hfff00113;
        ram_cell[    1164] = 32'h00209463;
        ram_cell[    1165] = 32'h0940106f;
        ram_cell[    1166] = 32'h00120213;
        ram_cell[    1167] = 32'h00200293;
        ram_cell[    1168] = 32'hfe5212e3;
        ram_cell[    1169] = 32'h07900193;
        ram_cell[    1170] = 32'h00000213;
        ram_cell[    1171] = 32'h00000093;
        ram_cell[    1172] = 32'h00000013;
        ram_cell[    1173] = 32'hfff00113;
        ram_cell[    1174] = 32'h00000013;
        ram_cell[    1175] = 32'h00209463;
        ram_cell[    1176] = 32'h0680106f;
        ram_cell[    1177] = 32'h00120213;
        ram_cell[    1178] = 32'h00200293;
        ram_cell[    1179] = 32'hfe5210e3;
        ram_cell[    1180] = 32'h07a00193;
        ram_cell[    1181] = 32'h00000213;
        ram_cell[    1182] = 32'h00000093;
        ram_cell[    1183] = 32'h00000013;
        ram_cell[    1184] = 32'h00000013;
        ram_cell[    1185] = 32'hfff00113;
        ram_cell[    1186] = 32'h00209463;
        ram_cell[    1187] = 32'h03c0106f;
        ram_cell[    1188] = 32'h00120213;
        ram_cell[    1189] = 32'h00200293;
        ram_cell[    1190] = 32'hfe5210e3;
        ram_cell[    1191] = 32'h00100093;
        ram_cell[    1192] = 32'h00000a63;
        ram_cell[    1193] = 32'h00108093;
        ram_cell[    1194] = 32'h00108093;
        ram_cell[    1195] = 32'h00108093;
        ram_cell[    1196] = 32'h00108093;
        ram_cell[    1197] = 32'h00108093;
        ram_cell[    1198] = 32'h00108093;
        ram_cell[    1199] = 32'h00300e93;
        ram_cell[    1200] = 32'h07b00193;
        ram_cell[    1201] = 32'h01d08463;
        ram_cell[    1202] = 32'h0000106f;
        ram_cell[    1203] = 32'h07c00193;
        ram_cell[    1204] = 32'h00000093;
        ram_cell[    1205] = 32'h00000113;
        ram_cell[    1206] = 32'h0020d663;
        ram_cell[    1207] = 32'h7e3016e3;
        ram_cell[    1208] = 32'h00301663;
        ram_cell[    1209] = 32'hfe20dee3;
        ram_cell[    1210] = 32'h7e3010e3;
        ram_cell[    1211] = 32'h07d00193;
        ram_cell[    1212] = 32'h00100093;
        ram_cell[    1213] = 32'h00100113;
        ram_cell[    1214] = 32'h0020d663;
        ram_cell[    1215] = 32'h7c3016e3;
        ram_cell[    1216] = 32'h00301663;
        ram_cell[    1217] = 32'hfe20dee3;
        ram_cell[    1218] = 32'h7c3010e3;
        ram_cell[    1219] = 32'h07e00193;
        ram_cell[    1220] = 32'hfff00093;
        ram_cell[    1221] = 32'hfff00113;
        ram_cell[    1222] = 32'h0020d663;
        ram_cell[    1223] = 32'h7a3016e3;
        ram_cell[    1224] = 32'h00301663;
        ram_cell[    1225] = 32'hfe20dee3;
        ram_cell[    1226] = 32'h7a3010e3;
        ram_cell[    1227] = 32'h07f00193;
        ram_cell[    1228] = 32'h00100093;
        ram_cell[    1229] = 32'h00000113;
        ram_cell[    1230] = 32'h0020d663;
        ram_cell[    1231] = 32'h783016e3;
        ram_cell[    1232] = 32'h00301663;
        ram_cell[    1233] = 32'hfe20dee3;
        ram_cell[    1234] = 32'h783010e3;
        ram_cell[    1235] = 32'h08000193;
        ram_cell[    1236] = 32'h00100093;
        ram_cell[    1237] = 32'hfff00113;
        ram_cell[    1238] = 32'h0020d663;
        ram_cell[    1239] = 32'h763016e3;
        ram_cell[    1240] = 32'h00301663;
        ram_cell[    1241] = 32'hfe20dee3;
        ram_cell[    1242] = 32'h763010e3;
        ram_cell[    1243] = 32'h08100193;
        ram_cell[    1244] = 32'hfff00093;
        ram_cell[    1245] = 32'hffe00113;
        ram_cell[    1246] = 32'h0020d663;
        ram_cell[    1247] = 32'h743016e3;
        ram_cell[    1248] = 32'h00301663;
        ram_cell[    1249] = 32'hfe20dee3;
        ram_cell[    1250] = 32'h743010e3;
        ram_cell[    1251] = 32'h08200193;
        ram_cell[    1252] = 32'h00000093;
        ram_cell[    1253] = 32'h00100113;
        ram_cell[    1254] = 32'h0020d463;
        ram_cell[    1255] = 32'h00301463;
        ram_cell[    1256] = 32'h723014e3;
        ram_cell[    1257] = 32'hfe20dee3;
        ram_cell[    1258] = 32'h08300193;
        ram_cell[    1259] = 32'hfff00093;
        ram_cell[    1260] = 32'h00100113;
        ram_cell[    1261] = 32'h0020d463;
        ram_cell[    1262] = 32'h00301463;
        ram_cell[    1263] = 32'h703016e3;
        ram_cell[    1264] = 32'hfe20dee3;
        ram_cell[    1265] = 32'h08400193;
        ram_cell[    1266] = 32'hffe00093;
        ram_cell[    1267] = 32'hfff00113;
        ram_cell[    1268] = 32'h0020d463;
        ram_cell[    1269] = 32'h00301463;
        ram_cell[    1270] = 32'h6e3018e3;
        ram_cell[    1271] = 32'hfe20dee3;
        ram_cell[    1272] = 32'h08500193;
        ram_cell[    1273] = 32'hffe00093;
        ram_cell[    1274] = 32'h00100113;
        ram_cell[    1275] = 32'h0020d463;
        ram_cell[    1276] = 32'h00301463;
        ram_cell[    1277] = 32'h6c301ae3;
        ram_cell[    1278] = 32'hfe20dee3;
        ram_cell[    1279] = 32'h08600193;
        ram_cell[    1280] = 32'h00000213;
        ram_cell[    1281] = 32'hfff00093;
        ram_cell[    1282] = 32'h00000113;
        ram_cell[    1283] = 32'h6a20dee3;
        ram_cell[    1284] = 32'h00120213;
        ram_cell[    1285] = 32'h00200293;
        ram_cell[    1286] = 32'hfe5216e3;
        ram_cell[    1287] = 32'h08700193;
        ram_cell[    1288] = 32'h00000213;
        ram_cell[    1289] = 32'hfff00093;
        ram_cell[    1290] = 32'h00000113;
        ram_cell[    1291] = 32'h00000013;
        ram_cell[    1292] = 32'h6820dce3;
        ram_cell[    1293] = 32'h00120213;
        ram_cell[    1294] = 32'h00200293;
        ram_cell[    1295] = 32'hfe5214e3;
        ram_cell[    1296] = 32'h08800193;
        ram_cell[    1297] = 32'h00000213;
        ram_cell[    1298] = 32'hfff00093;
        ram_cell[    1299] = 32'h00000113;
        ram_cell[    1300] = 32'h00000013;
        ram_cell[    1301] = 32'h00000013;
        ram_cell[    1302] = 32'h6620d8e3;
        ram_cell[    1303] = 32'h00120213;
        ram_cell[    1304] = 32'h00200293;
        ram_cell[    1305] = 32'hfe5212e3;
        ram_cell[    1306] = 32'h08900193;
        ram_cell[    1307] = 32'h00000213;
        ram_cell[    1308] = 32'hfff00093;
        ram_cell[    1309] = 32'h00000013;
        ram_cell[    1310] = 32'h00000113;
        ram_cell[    1311] = 32'h6420d6e3;
        ram_cell[    1312] = 32'h00120213;
        ram_cell[    1313] = 32'h00200293;
        ram_cell[    1314] = 32'hfe5214e3;
        ram_cell[    1315] = 32'h08a00193;
        ram_cell[    1316] = 32'h00000213;
        ram_cell[    1317] = 32'hfff00093;
        ram_cell[    1318] = 32'h00000013;
        ram_cell[    1319] = 32'h00000113;
        ram_cell[    1320] = 32'h00000013;
        ram_cell[    1321] = 32'h6220d2e3;
        ram_cell[    1322] = 32'h00120213;
        ram_cell[    1323] = 32'h00200293;
        ram_cell[    1324] = 32'hfe5212e3;
        ram_cell[    1325] = 32'h08b00193;
        ram_cell[    1326] = 32'h00000213;
        ram_cell[    1327] = 32'hfff00093;
        ram_cell[    1328] = 32'h00000013;
        ram_cell[    1329] = 32'h00000013;
        ram_cell[    1330] = 32'h00000113;
        ram_cell[    1331] = 32'h5e20dee3;
        ram_cell[    1332] = 32'h00120213;
        ram_cell[    1333] = 32'h00200293;
        ram_cell[    1334] = 32'hfe5212e3;
        ram_cell[    1335] = 32'h08c00193;
        ram_cell[    1336] = 32'h00000213;
        ram_cell[    1337] = 32'hfff00093;
        ram_cell[    1338] = 32'h00000113;
        ram_cell[    1339] = 32'h5c20dee3;
        ram_cell[    1340] = 32'h00120213;
        ram_cell[    1341] = 32'h00200293;
        ram_cell[    1342] = 32'hfe5216e3;
        ram_cell[    1343] = 32'h08d00193;
        ram_cell[    1344] = 32'h00000213;
        ram_cell[    1345] = 32'hfff00093;
        ram_cell[    1346] = 32'h00000113;
        ram_cell[    1347] = 32'h00000013;
        ram_cell[    1348] = 32'h5a20dce3;
        ram_cell[    1349] = 32'h00120213;
        ram_cell[    1350] = 32'h00200293;
        ram_cell[    1351] = 32'hfe5214e3;
        ram_cell[    1352] = 32'h08e00193;
        ram_cell[    1353] = 32'h00000213;
        ram_cell[    1354] = 32'hfff00093;
        ram_cell[    1355] = 32'h00000113;
        ram_cell[    1356] = 32'h00000013;
        ram_cell[    1357] = 32'h00000013;
        ram_cell[    1358] = 32'h5820d8e3;
        ram_cell[    1359] = 32'h00120213;
        ram_cell[    1360] = 32'h00200293;
        ram_cell[    1361] = 32'hfe5212e3;
        ram_cell[    1362] = 32'h08f00193;
        ram_cell[    1363] = 32'h00000213;
        ram_cell[    1364] = 32'hfff00093;
        ram_cell[    1365] = 32'h00000013;
        ram_cell[    1366] = 32'h00000113;
        ram_cell[    1367] = 32'h5620d6e3;
        ram_cell[    1368] = 32'h00120213;
        ram_cell[    1369] = 32'h00200293;
        ram_cell[    1370] = 32'hfe5214e3;
        ram_cell[    1371] = 32'h09000193;
        ram_cell[    1372] = 32'h00000213;
        ram_cell[    1373] = 32'hfff00093;
        ram_cell[    1374] = 32'h00000013;
        ram_cell[    1375] = 32'h00000113;
        ram_cell[    1376] = 32'h00000013;
        ram_cell[    1377] = 32'h5420d2e3;
        ram_cell[    1378] = 32'h00120213;
        ram_cell[    1379] = 32'h00200293;
        ram_cell[    1380] = 32'hfe5212e3;
        ram_cell[    1381] = 32'h09100193;
        ram_cell[    1382] = 32'h00000213;
        ram_cell[    1383] = 32'hfff00093;
        ram_cell[    1384] = 32'h00000013;
        ram_cell[    1385] = 32'h00000013;
        ram_cell[    1386] = 32'h00000113;
        ram_cell[    1387] = 32'h5020dee3;
        ram_cell[    1388] = 32'h00120213;
        ram_cell[    1389] = 32'h00200293;
        ram_cell[    1390] = 32'hfe5212e3;
        ram_cell[    1391] = 32'h00100093;
        ram_cell[    1392] = 32'h0000da63;
        ram_cell[    1393] = 32'h00108093;
        ram_cell[    1394] = 32'h00108093;
        ram_cell[    1395] = 32'h00108093;
        ram_cell[    1396] = 32'h00108093;
        ram_cell[    1397] = 32'h00108093;
        ram_cell[    1398] = 32'h00108093;
        ram_cell[    1399] = 32'h00300e93;
        ram_cell[    1400] = 32'h09200193;
        ram_cell[    1401] = 32'h4fd092e3;
        ram_cell[    1402] = 32'h09300193;
        ram_cell[    1403] = 32'h00000093;
        ram_cell[    1404] = 32'h00000113;
        ram_cell[    1405] = 32'h0020f663;
        ram_cell[    1406] = 32'h4c3018e3;
        ram_cell[    1407] = 32'h00301663;
        ram_cell[    1408] = 32'hfe20fee3;
        ram_cell[    1409] = 32'h4c3012e3;
        ram_cell[    1410] = 32'h09400193;
        ram_cell[    1411] = 32'h00100093;
        ram_cell[    1412] = 32'h00100113;
        ram_cell[    1413] = 32'h0020f663;
        ram_cell[    1414] = 32'h4a3018e3;
        ram_cell[    1415] = 32'h00301663;
        ram_cell[    1416] = 32'hfe20fee3;
        ram_cell[    1417] = 32'h4a3012e3;
        ram_cell[    1418] = 32'h09500193;
        ram_cell[    1419] = 32'hfff00093;
        ram_cell[    1420] = 32'hfff00113;
        ram_cell[    1421] = 32'h0020f663;
        ram_cell[    1422] = 32'h483018e3;
        ram_cell[    1423] = 32'h00301663;
        ram_cell[    1424] = 32'hfe20fee3;
        ram_cell[    1425] = 32'h483012e3;
        ram_cell[    1426] = 32'h09600193;
        ram_cell[    1427] = 32'h00100093;
        ram_cell[    1428] = 32'h00000113;
        ram_cell[    1429] = 32'h0020f663;
        ram_cell[    1430] = 32'h463018e3;
        ram_cell[    1431] = 32'h00301663;
        ram_cell[    1432] = 32'hfe20fee3;
        ram_cell[    1433] = 32'h463012e3;
        ram_cell[    1434] = 32'h09700193;
        ram_cell[    1435] = 32'hfff00093;
        ram_cell[    1436] = 32'hffe00113;
        ram_cell[    1437] = 32'h0020f663;
        ram_cell[    1438] = 32'h443018e3;
        ram_cell[    1439] = 32'h00301663;
        ram_cell[    1440] = 32'hfe20fee3;
        ram_cell[    1441] = 32'h443012e3;
        ram_cell[    1442] = 32'h09800193;
        ram_cell[    1443] = 32'hfff00093;
        ram_cell[    1444] = 32'h00000113;
        ram_cell[    1445] = 32'h0020f663;
        ram_cell[    1446] = 32'h423018e3;
        ram_cell[    1447] = 32'h00301663;
        ram_cell[    1448] = 32'hfe20fee3;
        ram_cell[    1449] = 32'h423012e3;
        ram_cell[    1450] = 32'h09900193;
        ram_cell[    1451] = 32'h00000093;
        ram_cell[    1452] = 32'h00100113;
        ram_cell[    1453] = 32'h0020f463;
        ram_cell[    1454] = 32'h00301463;
        ram_cell[    1455] = 32'h403016e3;
        ram_cell[    1456] = 32'hfe20fee3;
        ram_cell[    1457] = 32'h09a00193;
        ram_cell[    1458] = 32'hffe00093;
        ram_cell[    1459] = 32'hfff00113;
        ram_cell[    1460] = 32'h0020f463;
        ram_cell[    1461] = 32'h00301463;
        ram_cell[    1462] = 32'h3e3018e3;
        ram_cell[    1463] = 32'hfe20fee3;
        ram_cell[    1464] = 32'h09b00193;
        ram_cell[    1465] = 32'h00000093;
        ram_cell[    1466] = 32'hfff00113;
        ram_cell[    1467] = 32'h0020f463;
        ram_cell[    1468] = 32'h00301463;
        ram_cell[    1469] = 32'h3c301ae3;
        ram_cell[    1470] = 32'hfe20fee3;
        ram_cell[    1471] = 32'h09c00193;
        ram_cell[    1472] = 32'h800000b7;
        ram_cell[    1473] = 32'hfff08093;
        ram_cell[    1474] = 32'h80000137;
        ram_cell[    1475] = 32'h0020f463;
        ram_cell[    1476] = 32'h00301463;
        ram_cell[    1477] = 32'h3a301ae3;
        ram_cell[    1478] = 32'hfe20fee3;
        ram_cell[    1479] = 32'h09d00193;
        ram_cell[    1480] = 32'h00000213;
        ram_cell[    1481] = 32'hf00000b7;
        ram_cell[    1482] = 32'hfff08093;
        ram_cell[    1483] = 32'hf0000137;
        ram_cell[    1484] = 32'h3820fce3;
        ram_cell[    1485] = 32'h00120213;
        ram_cell[    1486] = 32'h00200293;
        ram_cell[    1487] = 32'hfe5214e3;
        ram_cell[    1488] = 32'h09e00193;
        ram_cell[    1489] = 32'h00000213;
        ram_cell[    1490] = 32'hf00000b7;
        ram_cell[    1491] = 32'hfff08093;
        ram_cell[    1492] = 32'hf0000137;
        ram_cell[    1493] = 32'h00000013;
        ram_cell[    1494] = 32'h3620f8e3;
        ram_cell[    1495] = 32'h00120213;
        ram_cell[    1496] = 32'h00200293;
        ram_cell[    1497] = 32'hfe5212e3;
        ram_cell[    1498] = 32'h09f00193;
        ram_cell[    1499] = 32'h00000213;
        ram_cell[    1500] = 32'hf00000b7;
        ram_cell[    1501] = 32'hfff08093;
        ram_cell[    1502] = 32'hf0000137;
        ram_cell[    1503] = 32'h00000013;
        ram_cell[    1504] = 32'h00000013;
        ram_cell[    1505] = 32'h3420f2e3;
        ram_cell[    1506] = 32'h00120213;
        ram_cell[    1507] = 32'h00200293;
        ram_cell[    1508] = 32'hfe5210e3;
        ram_cell[    1509] = 32'h0a000193;
        ram_cell[    1510] = 32'h00000213;
        ram_cell[    1511] = 32'hf00000b7;
        ram_cell[    1512] = 32'hfff08093;
        ram_cell[    1513] = 32'h00000013;
        ram_cell[    1514] = 32'hf0000137;
        ram_cell[    1515] = 32'h3020fee3;
        ram_cell[    1516] = 32'h00120213;
        ram_cell[    1517] = 32'h00200293;
        ram_cell[    1518] = 32'hfe5212e3;
        ram_cell[    1519] = 32'h0a100193;
        ram_cell[    1520] = 32'h00000213;
        ram_cell[    1521] = 32'hf00000b7;
        ram_cell[    1522] = 32'hfff08093;
        ram_cell[    1523] = 32'h00000013;
        ram_cell[    1524] = 32'hf0000137;
        ram_cell[    1525] = 32'h00000013;
        ram_cell[    1526] = 32'h2e20f8e3;
        ram_cell[    1527] = 32'h00120213;
        ram_cell[    1528] = 32'h00200293;
        ram_cell[    1529] = 32'hfe5210e3;
        ram_cell[    1530] = 32'h0a200193;
        ram_cell[    1531] = 32'h00000213;
        ram_cell[    1532] = 32'hf00000b7;
        ram_cell[    1533] = 32'hfff08093;
        ram_cell[    1534] = 32'h00000013;
        ram_cell[    1535] = 32'h00000013;
        ram_cell[    1536] = 32'hf0000137;
        ram_cell[    1537] = 32'h2c20f2e3;
        ram_cell[    1538] = 32'h00120213;
        ram_cell[    1539] = 32'h00200293;
        ram_cell[    1540] = 32'hfe5210e3;
        ram_cell[    1541] = 32'h0a300193;
        ram_cell[    1542] = 32'h00000213;
        ram_cell[    1543] = 32'hf00000b7;
        ram_cell[    1544] = 32'hfff08093;
        ram_cell[    1545] = 32'hf0000137;
        ram_cell[    1546] = 32'h2a20f0e3;
        ram_cell[    1547] = 32'h00120213;
        ram_cell[    1548] = 32'h00200293;
        ram_cell[    1549] = 32'hfe5214e3;
        ram_cell[    1550] = 32'h0a400193;
        ram_cell[    1551] = 32'h00000213;
        ram_cell[    1552] = 32'hf00000b7;
        ram_cell[    1553] = 32'hfff08093;
        ram_cell[    1554] = 32'hf0000137;
        ram_cell[    1555] = 32'h00000013;
        ram_cell[    1556] = 32'h2620fce3;
        ram_cell[    1557] = 32'h00120213;
        ram_cell[    1558] = 32'h00200293;
        ram_cell[    1559] = 32'hfe5212e3;
        ram_cell[    1560] = 32'h0a500193;
        ram_cell[    1561] = 32'h00000213;
        ram_cell[    1562] = 32'hf00000b7;
        ram_cell[    1563] = 32'hfff08093;
        ram_cell[    1564] = 32'hf0000137;
        ram_cell[    1565] = 32'h00000013;
        ram_cell[    1566] = 32'h00000013;
        ram_cell[    1567] = 32'h2420f6e3;
        ram_cell[    1568] = 32'h00120213;
        ram_cell[    1569] = 32'h00200293;
        ram_cell[    1570] = 32'hfe5210e3;
        ram_cell[    1571] = 32'h0a600193;
        ram_cell[    1572] = 32'h00000213;
        ram_cell[    1573] = 32'hf00000b7;
        ram_cell[    1574] = 32'hfff08093;
        ram_cell[    1575] = 32'h00000013;
        ram_cell[    1576] = 32'hf0000137;
        ram_cell[    1577] = 32'h2220f2e3;
        ram_cell[    1578] = 32'h00120213;
        ram_cell[    1579] = 32'h00200293;
        ram_cell[    1580] = 32'hfe5212e3;
        ram_cell[    1581] = 32'h0a700193;
        ram_cell[    1582] = 32'h00000213;
        ram_cell[    1583] = 32'hf00000b7;
        ram_cell[    1584] = 32'hfff08093;
        ram_cell[    1585] = 32'h00000013;
        ram_cell[    1586] = 32'hf0000137;
        ram_cell[    1587] = 32'h00000013;
        ram_cell[    1588] = 32'h1e20fce3;
        ram_cell[    1589] = 32'h00120213;
        ram_cell[    1590] = 32'h00200293;
        ram_cell[    1591] = 32'hfe5210e3;
        ram_cell[    1592] = 32'h0a800193;
        ram_cell[    1593] = 32'h00000213;
        ram_cell[    1594] = 32'hf00000b7;
        ram_cell[    1595] = 32'hfff08093;
        ram_cell[    1596] = 32'h00000013;
        ram_cell[    1597] = 32'h00000013;
        ram_cell[    1598] = 32'hf0000137;
        ram_cell[    1599] = 32'h1c20f6e3;
        ram_cell[    1600] = 32'h00120213;
        ram_cell[    1601] = 32'h00200293;
        ram_cell[    1602] = 32'hfe5210e3;
        ram_cell[    1603] = 32'h00100093;
        ram_cell[    1604] = 32'h0000fa63;
        ram_cell[    1605] = 32'h00108093;
        ram_cell[    1606] = 32'h00108093;
        ram_cell[    1607] = 32'h00108093;
        ram_cell[    1608] = 32'h00108093;
        ram_cell[    1609] = 32'h00108093;
        ram_cell[    1610] = 32'h00108093;
        ram_cell[    1611] = 32'h00300e93;
        ram_cell[    1612] = 32'h0a900193;
        ram_cell[    1613] = 32'h19d09ae3;
        ram_cell[    1614] = 32'h0aa00193;
        ram_cell[    1615] = 32'h00000093;
        ram_cell[    1616] = 32'h00100113;
        ram_cell[    1617] = 32'h0020c663;
        ram_cell[    1618] = 32'h183010e3;
        ram_cell[    1619] = 32'h00301663;
        ram_cell[    1620] = 32'hfe20cee3;
        ram_cell[    1621] = 32'h16301ae3;
        ram_cell[    1622] = 32'h0ab00193;
        ram_cell[    1623] = 32'hfff00093;
        ram_cell[    1624] = 32'h00100113;
        ram_cell[    1625] = 32'h0020c663;
        ram_cell[    1626] = 32'h163010e3;
        ram_cell[    1627] = 32'h00301663;
        ram_cell[    1628] = 32'hfe20cee3;
        ram_cell[    1629] = 32'h14301ae3;
        ram_cell[    1630] = 32'h0ac00193;
        ram_cell[    1631] = 32'hffe00093;
        ram_cell[    1632] = 32'hfff00113;
        ram_cell[    1633] = 32'h0020c663;
        ram_cell[    1634] = 32'h143010e3;
        ram_cell[    1635] = 32'h00301663;
        ram_cell[    1636] = 32'hfe20cee3;
        ram_cell[    1637] = 32'h12301ae3;
        ram_cell[    1638] = 32'h0ad00193;
        ram_cell[    1639] = 32'h00100093;
        ram_cell[    1640] = 32'h00000113;
        ram_cell[    1641] = 32'h0020c463;
        ram_cell[    1642] = 32'h00301463;
        ram_cell[    1643] = 32'h10301ee3;
        ram_cell[    1644] = 32'hfe20cee3;
        ram_cell[    1645] = 32'h0ae00193;
        ram_cell[    1646] = 32'h00100093;
        ram_cell[    1647] = 32'hfff00113;
        ram_cell[    1648] = 32'h0020c463;
        ram_cell[    1649] = 32'h00301463;
        ram_cell[    1650] = 32'h103010e3;
        ram_cell[    1651] = 32'hfe20cee3;
        ram_cell[    1652] = 32'h0af00193;
        ram_cell[    1653] = 32'hfff00093;
        ram_cell[    1654] = 32'hffe00113;
        ram_cell[    1655] = 32'h0020c463;
        ram_cell[    1656] = 32'h00301463;
        ram_cell[    1657] = 32'h0e3012e3;
        ram_cell[    1658] = 32'hfe20cee3;
        ram_cell[    1659] = 32'h0b000193;
        ram_cell[    1660] = 32'h00100093;
        ram_cell[    1661] = 32'hffe00113;
        ram_cell[    1662] = 32'h0020c463;
        ram_cell[    1663] = 32'h00301463;
        ram_cell[    1664] = 32'h0c3014e3;
        ram_cell[    1665] = 32'hfe20cee3;
        ram_cell[    1666] = 32'h0b100193;
        ram_cell[    1667] = 32'h00000213;
        ram_cell[    1668] = 32'h00000093;
        ram_cell[    1669] = 32'hfff00113;
        ram_cell[    1670] = 32'h0a20c8e3;
        ram_cell[    1671] = 32'h00120213;
        ram_cell[    1672] = 32'h00200293;
        ram_cell[    1673] = 32'hfe5216e3;
        ram_cell[    1674] = 32'h0b200193;
        ram_cell[    1675] = 32'h00000213;
        ram_cell[    1676] = 32'h00000093;
        ram_cell[    1677] = 32'hfff00113;
        ram_cell[    1678] = 32'h00000013;
        ram_cell[    1679] = 32'h0820c6e3;
        ram_cell[    1680] = 32'h00120213;
        ram_cell[    1681] = 32'h00200293;
        ram_cell[    1682] = 32'hfe5214e3;
        ram_cell[    1683] = 32'h0b300193;
        ram_cell[    1684] = 32'h00000213;
        ram_cell[    1685] = 32'h00000093;
        ram_cell[    1686] = 32'hfff00113;
        ram_cell[    1687] = 32'h00000013;
        ram_cell[    1688] = 32'h00000013;
        ram_cell[    1689] = 32'h0620c2e3;
        ram_cell[    1690] = 32'h00120213;
        ram_cell[    1691] = 32'h00200293;
        ram_cell[    1692] = 32'hfe5212e3;
        ram_cell[    1693] = 32'h0b400193;
        ram_cell[    1694] = 32'h00000213;
        ram_cell[    1695] = 32'h00000093;
        ram_cell[    1696] = 32'h00000013;
        ram_cell[    1697] = 32'hfff00113;
        ram_cell[    1698] = 32'h0420c0e3;
        ram_cell[    1699] = 32'h00120213;
        ram_cell[    1700] = 32'h00200293;
        ram_cell[    1701] = 32'hfe5214e3;
        ram_cell[    1702] = 32'h0b500193;
        ram_cell[    1703] = 32'h00000213;
        ram_cell[    1704] = 32'h00000093;
        ram_cell[    1705] = 32'h00000013;
        ram_cell[    1706] = 32'hfff00113;
        ram_cell[    1707] = 32'h00000013;
        ram_cell[    1708] = 32'h0020cce3;
        ram_cell[    1709] = 32'h00120213;
        ram_cell[    1710] = 32'h00200293;
        ram_cell[    1711] = 32'hfe5212e3;
        ram_cell[    1712] = 32'h0b600193;
        ram_cell[    1713] = 32'h00000213;
        ram_cell[    1714] = 32'h00000093;
        ram_cell[    1715] = 32'h00000013;
        ram_cell[    1716] = 32'h00000013;
        ram_cell[    1717] = 32'hfff00113;
        ram_cell[    1718] = 32'h7e20c863;
        ram_cell[    1719] = 32'h00120213;
        ram_cell[    1720] = 32'h00200293;
        ram_cell[    1721] = 32'hfe5212e3;
        ram_cell[    1722] = 32'h0b700193;
        ram_cell[    1723] = 32'h00000213;
        ram_cell[    1724] = 32'h00000093;
        ram_cell[    1725] = 32'hfff00113;
        ram_cell[    1726] = 32'h7c20c863;
        ram_cell[    1727] = 32'h00120213;
        ram_cell[    1728] = 32'h00200293;
        ram_cell[    1729] = 32'hfe5216e3;
        ram_cell[    1730] = 32'h0b800193;
        ram_cell[    1731] = 32'h00000213;
        ram_cell[    1732] = 32'h00000093;
        ram_cell[    1733] = 32'hfff00113;
        ram_cell[    1734] = 32'h00000013;
        ram_cell[    1735] = 32'h7a20c663;
        ram_cell[    1736] = 32'h00120213;
        ram_cell[    1737] = 32'h00200293;
        ram_cell[    1738] = 32'hfe5214e3;
        ram_cell[    1739] = 32'h0b900193;
        ram_cell[    1740] = 32'h00000213;
        ram_cell[    1741] = 32'h00000093;
        ram_cell[    1742] = 32'hfff00113;
        ram_cell[    1743] = 32'h00000013;
        ram_cell[    1744] = 32'h00000013;
        ram_cell[    1745] = 32'h7820c263;
        ram_cell[    1746] = 32'h00120213;
        ram_cell[    1747] = 32'h00200293;
        ram_cell[    1748] = 32'hfe5212e3;
        ram_cell[    1749] = 32'h0ba00193;
        ram_cell[    1750] = 32'h00000213;
        ram_cell[    1751] = 32'h00000093;
        ram_cell[    1752] = 32'h00000013;
        ram_cell[    1753] = 32'hfff00113;
        ram_cell[    1754] = 32'h7620c063;
        ram_cell[    1755] = 32'h00120213;
        ram_cell[    1756] = 32'h00200293;
        ram_cell[    1757] = 32'hfe5214e3;
        ram_cell[    1758] = 32'h0bb00193;
        ram_cell[    1759] = 32'h00000213;
        ram_cell[    1760] = 32'h00000093;
        ram_cell[    1761] = 32'h00000013;
        ram_cell[    1762] = 32'hfff00113;
        ram_cell[    1763] = 32'h00000013;
        ram_cell[    1764] = 32'h7220cc63;
        ram_cell[    1765] = 32'h00120213;
        ram_cell[    1766] = 32'h00200293;
        ram_cell[    1767] = 32'hfe5212e3;
        ram_cell[    1768] = 32'h0bc00193;
        ram_cell[    1769] = 32'h00000213;
        ram_cell[    1770] = 32'h00000093;
        ram_cell[    1771] = 32'h00000013;
        ram_cell[    1772] = 32'h00000013;
        ram_cell[    1773] = 32'hfff00113;
        ram_cell[    1774] = 32'h7020c863;
        ram_cell[    1775] = 32'h00120213;
        ram_cell[    1776] = 32'h00200293;
        ram_cell[    1777] = 32'hfe5212e3;
        ram_cell[    1778] = 32'h00100093;
        ram_cell[    1779] = 32'h00104a63;
        ram_cell[    1780] = 32'h00108093;
        ram_cell[    1781] = 32'h00108093;
        ram_cell[    1782] = 32'h00108093;
        ram_cell[    1783] = 32'h00108093;
        ram_cell[    1784] = 32'h00108093;
        ram_cell[    1785] = 32'h00108093;
        ram_cell[    1786] = 32'h00300e93;
        ram_cell[    1787] = 32'h0bd00193;
        ram_cell[    1788] = 32'h6dd09c63;
        ram_cell[    1789] = 32'h0be00193;
        ram_cell[    1790] = 32'h00000093;
        ram_cell[    1791] = 32'h00100113;
        ram_cell[    1792] = 32'h0020e663;
        ram_cell[    1793] = 32'h6c301263;
        ram_cell[    1794] = 32'h00301663;
        ram_cell[    1795] = 32'hfe20eee3;
        ram_cell[    1796] = 32'h6a301c63;
        ram_cell[    1797] = 32'h0bf00193;
        ram_cell[    1798] = 32'hffe00093;
        ram_cell[    1799] = 32'hfff00113;
        ram_cell[    1800] = 32'h0020e663;
        ram_cell[    1801] = 32'h6a301263;
        ram_cell[    1802] = 32'h00301663;
        ram_cell[    1803] = 32'hfe20eee3;
        ram_cell[    1804] = 32'h68301c63;
        ram_cell[    1805] = 32'h0c000193;
        ram_cell[    1806] = 32'h00000093;
        ram_cell[    1807] = 32'hfff00113;
        ram_cell[    1808] = 32'h0020e663;
        ram_cell[    1809] = 32'h68301263;
        ram_cell[    1810] = 32'h00301663;
        ram_cell[    1811] = 32'hfe20eee3;
        ram_cell[    1812] = 32'h66301c63;
        ram_cell[    1813] = 32'h0c100193;
        ram_cell[    1814] = 32'h00100093;
        ram_cell[    1815] = 32'h00000113;
        ram_cell[    1816] = 32'h0020e463;
        ram_cell[    1817] = 32'h00301463;
        ram_cell[    1818] = 32'h66301063;
        ram_cell[    1819] = 32'hfe20eee3;
        ram_cell[    1820] = 32'h0c200193;
        ram_cell[    1821] = 32'hfff00093;
        ram_cell[    1822] = 32'hffe00113;
        ram_cell[    1823] = 32'h0020e463;
        ram_cell[    1824] = 32'h00301463;
        ram_cell[    1825] = 32'h64301263;
        ram_cell[    1826] = 32'hfe20eee3;
        ram_cell[    1827] = 32'h0c300193;
        ram_cell[    1828] = 32'hfff00093;
        ram_cell[    1829] = 32'h00000113;
        ram_cell[    1830] = 32'h0020e463;
        ram_cell[    1831] = 32'h00301463;
        ram_cell[    1832] = 32'h62301463;
        ram_cell[    1833] = 32'hfe20eee3;
        ram_cell[    1834] = 32'h0c400193;
        ram_cell[    1835] = 32'h800000b7;
        ram_cell[    1836] = 32'h80000137;
        ram_cell[    1837] = 32'hfff10113;
        ram_cell[    1838] = 32'h0020e463;
        ram_cell[    1839] = 32'h00301463;
        ram_cell[    1840] = 32'h60301463;
        ram_cell[    1841] = 32'hfe20eee3;
        ram_cell[    1842] = 32'h0c500193;
        ram_cell[    1843] = 32'h00000213;
        ram_cell[    1844] = 32'hf00000b7;
        ram_cell[    1845] = 32'hf0000137;
        ram_cell[    1846] = 32'hfff10113;
        ram_cell[    1847] = 32'h5e20e663;
        ram_cell[    1848] = 32'h00120213;
        ram_cell[    1849] = 32'h00200293;
        ram_cell[    1850] = 32'hfe5214e3;
        ram_cell[    1851] = 32'h0c600193;
        ram_cell[    1852] = 32'h00000213;
        ram_cell[    1853] = 32'hf00000b7;
        ram_cell[    1854] = 32'hf0000137;
        ram_cell[    1855] = 32'hfff10113;
        ram_cell[    1856] = 32'h00000013;
        ram_cell[    1857] = 32'h5c20e263;
        ram_cell[    1858] = 32'h00120213;
        ram_cell[    1859] = 32'h00200293;
        ram_cell[    1860] = 32'hfe5212e3;
        ram_cell[    1861] = 32'h0c700193;
        ram_cell[    1862] = 32'h00000213;
        ram_cell[    1863] = 32'hf00000b7;
        ram_cell[    1864] = 32'hf0000137;
        ram_cell[    1865] = 32'hfff10113;
        ram_cell[    1866] = 32'h00000013;
        ram_cell[    1867] = 32'h00000013;
        ram_cell[    1868] = 32'h5820ec63;
        ram_cell[    1869] = 32'h00120213;
        ram_cell[    1870] = 32'h00200293;
        ram_cell[    1871] = 32'hfe5210e3;
        ram_cell[    1872] = 32'h0c800193;
        ram_cell[    1873] = 32'h00000213;
        ram_cell[    1874] = 32'hf00000b7;
        ram_cell[    1875] = 32'h00000013;
        ram_cell[    1876] = 32'hf0000137;
        ram_cell[    1877] = 32'hfff10113;
        ram_cell[    1878] = 32'h5620e863;
        ram_cell[    1879] = 32'h00120213;
        ram_cell[    1880] = 32'h00200293;
        ram_cell[    1881] = 32'hfe5212e3;
        ram_cell[    1882] = 32'h0c900193;
        ram_cell[    1883] = 32'h00000213;
        ram_cell[    1884] = 32'hf00000b7;
        ram_cell[    1885] = 32'h00000013;
        ram_cell[    1886] = 32'hf0000137;
        ram_cell[    1887] = 32'hfff10113;
        ram_cell[    1888] = 32'h00000013;
        ram_cell[    1889] = 32'h5420e263;
        ram_cell[    1890] = 32'h00120213;
        ram_cell[    1891] = 32'h00200293;
        ram_cell[    1892] = 32'hfe5210e3;
        ram_cell[    1893] = 32'h0ca00193;
        ram_cell[    1894] = 32'h00000213;
        ram_cell[    1895] = 32'hf00000b7;
        ram_cell[    1896] = 32'h00000013;
        ram_cell[    1897] = 32'h00000013;
        ram_cell[    1898] = 32'hf0000137;
        ram_cell[    1899] = 32'hfff10113;
        ram_cell[    1900] = 32'h5020ec63;
        ram_cell[    1901] = 32'h00120213;
        ram_cell[    1902] = 32'h00200293;
        ram_cell[    1903] = 32'hfe5210e3;
        ram_cell[    1904] = 32'h0cb00193;
        ram_cell[    1905] = 32'h00000213;
        ram_cell[    1906] = 32'hf00000b7;
        ram_cell[    1907] = 32'hf0000137;
        ram_cell[    1908] = 32'hfff10113;
        ram_cell[    1909] = 32'h4e20ea63;
        ram_cell[    1910] = 32'h00120213;
        ram_cell[    1911] = 32'h00200293;
        ram_cell[    1912] = 32'hfe5214e3;
        ram_cell[    1913] = 32'h0cc00193;
        ram_cell[    1914] = 32'h00000213;
        ram_cell[    1915] = 32'hf00000b7;
        ram_cell[    1916] = 32'hf0000137;
        ram_cell[    1917] = 32'hfff10113;
        ram_cell[    1918] = 32'h00000013;
        ram_cell[    1919] = 32'h4c20e663;
        ram_cell[    1920] = 32'h00120213;
        ram_cell[    1921] = 32'h00200293;
        ram_cell[    1922] = 32'hfe5212e3;
        ram_cell[    1923] = 32'h0cd00193;
        ram_cell[    1924] = 32'h00000213;
        ram_cell[    1925] = 32'hf00000b7;
        ram_cell[    1926] = 32'hf0000137;
        ram_cell[    1927] = 32'hfff10113;
        ram_cell[    1928] = 32'h00000013;
        ram_cell[    1929] = 32'h00000013;
        ram_cell[    1930] = 32'h4a20e063;
        ram_cell[    1931] = 32'h00120213;
        ram_cell[    1932] = 32'h00200293;
        ram_cell[    1933] = 32'hfe5210e3;
        ram_cell[    1934] = 32'h0ce00193;
        ram_cell[    1935] = 32'h00000213;
        ram_cell[    1936] = 32'hf00000b7;
        ram_cell[    1937] = 32'h00000013;
        ram_cell[    1938] = 32'hf0000137;
        ram_cell[    1939] = 32'hfff10113;
        ram_cell[    1940] = 32'h4620ec63;
        ram_cell[    1941] = 32'h00120213;
        ram_cell[    1942] = 32'h00200293;
        ram_cell[    1943] = 32'hfe5212e3;
        ram_cell[    1944] = 32'h0cf00193;
        ram_cell[    1945] = 32'h00000213;
        ram_cell[    1946] = 32'hf00000b7;
        ram_cell[    1947] = 32'h00000013;
        ram_cell[    1948] = 32'hf0000137;
        ram_cell[    1949] = 32'hfff10113;
        ram_cell[    1950] = 32'h00000013;
        ram_cell[    1951] = 32'h4420e663;
        ram_cell[    1952] = 32'h00120213;
        ram_cell[    1953] = 32'h00200293;
        ram_cell[    1954] = 32'hfe5210e3;
        ram_cell[    1955] = 32'h0d000193;
        ram_cell[    1956] = 32'h00000213;
        ram_cell[    1957] = 32'hf00000b7;
        ram_cell[    1958] = 32'h00000013;
        ram_cell[    1959] = 32'h00000013;
        ram_cell[    1960] = 32'hf0000137;
        ram_cell[    1961] = 32'hfff10113;
        ram_cell[    1962] = 32'h4220e063;
        ram_cell[    1963] = 32'h00120213;
        ram_cell[    1964] = 32'h00200293;
        ram_cell[    1965] = 32'hfe5210e3;
        ram_cell[    1966] = 32'h00100093;
        ram_cell[    1967] = 32'h00106a63;
        ram_cell[    1968] = 32'h00108093;
        ram_cell[    1969] = 32'h00108093;
        ram_cell[    1970] = 32'h00108093;
        ram_cell[    1971] = 32'h00108093;
        ram_cell[    1972] = 32'h00108093;
        ram_cell[    1973] = 32'h00108093;
        ram_cell[    1974] = 32'h00300e93;
        ram_cell[    1975] = 32'h0d100193;
        ram_cell[    1976] = 32'h3fd09463;
        ram_cell[    1977] = 32'h0d200193;
        ram_cell[    1978] = 32'h00000093;
        ram_cell[    1979] = 32'h00100113;
        ram_cell[    1980] = 32'h00209663;
        ram_cell[    1981] = 32'h3c301a63;
        ram_cell[    1982] = 32'h00301663;
        ram_cell[    1983] = 32'hfe209ee3;
        ram_cell[    1984] = 32'h3c301463;
        ram_cell[    1985] = 32'h0d300193;
        ram_cell[    1986] = 32'h00100093;
        ram_cell[    1987] = 32'h00000113;
        ram_cell[    1988] = 32'h00209663;
        ram_cell[    1989] = 32'h3a301a63;
        ram_cell[    1990] = 32'h00301663;
        ram_cell[    1991] = 32'hfe209ee3;
        ram_cell[    1992] = 32'h3a301463;
        ram_cell[    1993] = 32'h0d400193;
        ram_cell[    1994] = 32'hfff00093;
        ram_cell[    1995] = 32'h00100113;
        ram_cell[    1996] = 32'h00209663;
        ram_cell[    1997] = 32'h38301a63;
        ram_cell[    1998] = 32'h00301663;
        ram_cell[    1999] = 32'hfe209ee3;
        ram_cell[    2000] = 32'h38301463;
        ram_cell[    2001] = 32'h0d500193;
        ram_cell[    2002] = 32'h00100093;
        ram_cell[    2003] = 32'hfff00113;
        ram_cell[    2004] = 32'h00209663;
        ram_cell[    2005] = 32'h36301a63;
        ram_cell[    2006] = 32'h00301663;
        ram_cell[    2007] = 32'hfe209ee3;
        ram_cell[    2008] = 32'h36301463;
        ram_cell[    2009] = 32'h0d600193;
        ram_cell[    2010] = 32'h00000093;
        ram_cell[    2011] = 32'h00000113;
        ram_cell[    2012] = 32'h00209463;
        ram_cell[    2013] = 32'h00301463;
        ram_cell[    2014] = 32'h34301863;
        ram_cell[    2015] = 32'hfe209ee3;
        ram_cell[    2016] = 32'h0d700193;
        ram_cell[    2017] = 32'h00100093;
        ram_cell[    2018] = 32'h00100113;
        ram_cell[    2019] = 32'h00209463;
        ram_cell[    2020] = 32'h00301463;
        ram_cell[    2021] = 32'h32301a63;
        ram_cell[    2022] = 32'hfe209ee3;
        ram_cell[    2023] = 32'h0d800193;
        ram_cell[    2024] = 32'hfff00093;
        ram_cell[    2025] = 32'hfff00113;
        ram_cell[    2026] = 32'h00209463;
        ram_cell[    2027] = 32'h00301463;
        ram_cell[    2028] = 32'h30301c63;
        ram_cell[    2029] = 32'hfe209ee3;
        ram_cell[    2030] = 32'h0d900193;
        ram_cell[    2031] = 32'h00000213;
        ram_cell[    2032] = 32'h00000093;
        ram_cell[    2033] = 32'h00000113;
        ram_cell[    2034] = 32'h30209063;
        ram_cell[    2035] = 32'h00120213;
        ram_cell[    2036] = 32'h00200293;
        ram_cell[    2037] = 32'hfe5216e3;
        ram_cell[    2038] = 32'h0da00193;
        ram_cell[    2039] = 32'h00000213;
        ram_cell[    2040] = 32'h00000093;
        ram_cell[    2041] = 32'h00000113;
        ram_cell[    2042] = 32'h00000013;
        ram_cell[    2043] = 32'h2c209e63;
        ram_cell[    2044] = 32'h00120213;
        ram_cell[    2045] = 32'h00200293;
        ram_cell[    2046] = 32'hfe5214e3;
        ram_cell[    2047] = 32'h0db00193;
        ram_cell[    2048] = 32'h00000213;
        ram_cell[    2049] = 32'h00000093;
        ram_cell[    2050] = 32'h00000113;
        ram_cell[    2051] = 32'h00000013;
        ram_cell[    2052] = 32'h00000013;
        ram_cell[    2053] = 32'h2a209a63;
        ram_cell[    2054] = 32'h00120213;
        ram_cell[    2055] = 32'h00200293;
        ram_cell[    2056] = 32'hfe5212e3;
        ram_cell[    2057] = 32'h0dc00193;
        ram_cell[    2058] = 32'h00000213;
        ram_cell[    2059] = 32'h00000093;
        ram_cell[    2060] = 32'h00000013;
        ram_cell[    2061] = 32'h00000113;
        ram_cell[    2062] = 32'h28209863;
        ram_cell[    2063] = 32'h00120213;
        ram_cell[    2064] = 32'h00200293;
        ram_cell[    2065] = 32'hfe5214e3;
        ram_cell[    2066] = 32'h0dd00193;
        ram_cell[    2067] = 32'h00000213;
        ram_cell[    2068] = 32'h00000093;
        ram_cell[    2069] = 32'h00000013;
        ram_cell[    2070] = 32'h00000113;
        ram_cell[    2071] = 32'h00000013;
        ram_cell[    2072] = 32'h26209463;
        ram_cell[    2073] = 32'h00120213;
        ram_cell[    2074] = 32'h00200293;
        ram_cell[    2075] = 32'hfe5212e3;
        ram_cell[    2076] = 32'h0de00193;
        ram_cell[    2077] = 32'h00000213;
        ram_cell[    2078] = 32'h00000093;
        ram_cell[    2079] = 32'h00000013;
        ram_cell[    2080] = 32'h00000013;
        ram_cell[    2081] = 32'h00000113;
        ram_cell[    2082] = 32'h24209063;
        ram_cell[    2083] = 32'h00120213;
        ram_cell[    2084] = 32'h00200293;
        ram_cell[    2085] = 32'hfe5212e3;
        ram_cell[    2086] = 32'h0df00193;
        ram_cell[    2087] = 32'h00000213;
        ram_cell[    2088] = 32'h00000093;
        ram_cell[    2089] = 32'h00000113;
        ram_cell[    2090] = 32'h22209063;
        ram_cell[    2091] = 32'h00120213;
        ram_cell[    2092] = 32'h00200293;
        ram_cell[    2093] = 32'hfe5216e3;
        ram_cell[    2094] = 32'h0e000193;
        ram_cell[    2095] = 32'h00000213;
        ram_cell[    2096] = 32'h00000093;
        ram_cell[    2097] = 32'h00000113;
        ram_cell[    2098] = 32'h00000013;
        ram_cell[    2099] = 32'h1e209e63;
        ram_cell[    2100] = 32'h00120213;
        ram_cell[    2101] = 32'h00200293;
        ram_cell[    2102] = 32'hfe5214e3;
        ram_cell[    2103] = 32'h0e100193;
        ram_cell[    2104] = 32'h00000213;
        ram_cell[    2105] = 32'h00000093;
        ram_cell[    2106] = 32'h00000113;
        ram_cell[    2107] = 32'h00000013;
        ram_cell[    2108] = 32'h00000013;
        ram_cell[    2109] = 32'h1c209a63;
        ram_cell[    2110] = 32'h00120213;
        ram_cell[    2111] = 32'h00200293;
        ram_cell[    2112] = 32'hfe5212e3;
        ram_cell[    2113] = 32'h0e200193;
        ram_cell[    2114] = 32'h00000213;
        ram_cell[    2115] = 32'h00000093;
        ram_cell[    2116] = 32'h00000013;
        ram_cell[    2117] = 32'h00000113;
        ram_cell[    2118] = 32'h1a209863;
        ram_cell[    2119] = 32'h00120213;
        ram_cell[    2120] = 32'h00200293;
        ram_cell[    2121] = 32'hfe5214e3;
        ram_cell[    2122] = 32'h0e300193;
        ram_cell[    2123] = 32'h00000213;
        ram_cell[    2124] = 32'h00000093;
        ram_cell[    2125] = 32'h00000013;
        ram_cell[    2126] = 32'h00000113;
        ram_cell[    2127] = 32'h00000013;
        ram_cell[    2128] = 32'h18209463;
        ram_cell[    2129] = 32'h00120213;
        ram_cell[    2130] = 32'h00200293;
        ram_cell[    2131] = 32'hfe5212e3;
        ram_cell[    2132] = 32'h0e400193;
        ram_cell[    2133] = 32'h00000213;
        ram_cell[    2134] = 32'h00000093;
        ram_cell[    2135] = 32'h00000013;
        ram_cell[    2136] = 32'h00000013;
        ram_cell[    2137] = 32'h00000113;
        ram_cell[    2138] = 32'h16209063;
        ram_cell[    2139] = 32'h00120213;
        ram_cell[    2140] = 32'h00200293;
        ram_cell[    2141] = 32'hfe5212e3;
        ram_cell[    2142] = 32'h00100093;
        ram_cell[    2143] = 32'h00009a63;
        ram_cell[    2144] = 32'h00108093;
        ram_cell[    2145] = 32'h00108093;
        ram_cell[    2146] = 32'h00108093;
        ram_cell[    2147] = 32'h00108093;
        ram_cell[    2148] = 32'h00108093;
        ram_cell[    2149] = 32'h00108093;
        ram_cell[    2150] = 32'h00300e93;
        ram_cell[    2151] = 32'h0e500193;
        ram_cell[    2152] = 32'h13d09463;
        ram_cell[    2153] = 32'h00200193;
        ram_cell[    2154] = 32'h00000093;
        ram_cell[    2155] = 32'h0100026f;
        ram_cell[    2156] = 32'h00000013;
        ram_cell[    2157] = 32'h00000013;
        ram_cell[    2158] = 32'h1100006f;
        ram_cell[    2159] = 32'h00000317;
        ram_cell[    2160] = 32'hff430313;
        ram_cell[    2161] = 32'h10431263;
        ram_cell[    2162] = 32'h00100093;
        ram_cell[    2163] = 32'h0140006f;
        ram_cell[    2164] = 32'h00108093;
        ram_cell[    2165] = 32'h00108093;
        ram_cell[    2166] = 32'h00108093;
        ram_cell[    2167] = 32'h00108093;
        ram_cell[    2168] = 32'h00108093;
        ram_cell[    2169] = 32'h00108093;
        ram_cell[    2170] = 32'h00300e93;
        ram_cell[    2171] = 32'h0e800193;
        ram_cell[    2172] = 32'h0dd09c63;
        ram_cell[    2173] = 32'h00200193;
        ram_cell[    2174] = 32'h00000293;
        ram_cell[    2175] = 32'h00000317;
        ram_cell[    2176] = 32'h01030313;
        ram_cell[    2177] = 32'h000302e7;
        ram_cell[    2178] = 32'h0c00006f;
        ram_cell[    2179] = 32'h00000317;
        ram_cell[    2180] = 32'hffc30313;
        ram_cell[    2181] = 32'h0a629a63;
        ram_cell[    2182] = 32'h0e900193;
        ram_cell[    2183] = 32'h00000213;
        ram_cell[    2184] = 32'h00000317;
        ram_cell[    2185] = 32'h01030313;
        ram_cell[    2186] = 32'h000309e7;
        ram_cell[    2187] = 32'h08301e63;
        ram_cell[    2188] = 32'h00120213;
        ram_cell[    2189] = 32'h00200293;
        ram_cell[    2190] = 32'hfe5214e3;
        ram_cell[    2191] = 32'h0ea00193;
        ram_cell[    2192] = 32'h00000213;
        ram_cell[    2193] = 32'h00000317;
        ram_cell[    2194] = 32'h01430313;
        ram_cell[    2195] = 32'h00000013;
        ram_cell[    2196] = 32'h000309e7;
        ram_cell[    2197] = 32'h06301a63;
        ram_cell[    2198] = 32'h00120213;
        ram_cell[    2199] = 32'h00200293;
        ram_cell[    2200] = 32'hfe5212e3;
        ram_cell[    2201] = 32'h0eb00193;
        ram_cell[    2202] = 32'h00000213;
        ram_cell[    2203] = 32'h00000317;
        ram_cell[    2204] = 32'h01830313;
        ram_cell[    2205] = 32'h00000013;
        ram_cell[    2206] = 32'h00000013;
        ram_cell[    2207] = 32'h000309e7;
        ram_cell[    2208] = 32'h04301463;
        ram_cell[    2209] = 32'h00120213;
        ram_cell[    2210] = 32'h00200293;
        ram_cell[    2211] = 32'hfe5210e3;
        ram_cell[    2212] = 32'h00100293;
        ram_cell[    2213] = 32'h00000317;
        ram_cell[    2214] = 32'h01c30313;
        ram_cell[    2215] = 32'hffc30067;
        ram_cell[    2216] = 32'h00128293;
        ram_cell[    2217] = 32'h00128293;
        ram_cell[    2218] = 32'h00128293;
        ram_cell[    2219] = 32'h00128293;
        ram_cell[    2220] = 32'h00128293;
        ram_cell[    2221] = 32'h00128293;
        ram_cell[    2222] = 32'h00400e93;
        ram_cell[    2223] = 32'h0ec00193;
        ram_cell[    2224] = 32'h01d29463;
        ram_cell[    2225] = 32'h00301463;
        ram_cell[    2226] = 32'h00000a6f;
        ram_cell[    2227] = 32'h00100193;
        ram_cell[    2228] = 32'h00000a6f;
        ram_cell[    2229] = 32'hc0001073;
        ram_cell[    2230] = 32'h00000000;
        ram_cell[    2231] = 32'h00000000;
        ram_cell[    2232] = 32'h00000000;
        ram_cell[    2233] = 32'h00000000;
        ram_cell[    2234] = 32'h00000000;
        ram_cell[    2235] = 32'h00000000;
        ram_cell[    2236] = 32'h00000000;
        ram_cell[    2237] = 32'h00000000;
        ram_cell[    2238] = 32'h00000000;
        ram_cell[    2239] = 32'h00000000;
        ram_cell[    2240] = 32'h00000000;
        ram_cell[    2241] = 32'h00000000;
        ram_cell[    2242] = 32'h00000000;
        ram_cell[    2243] = 32'h00000000;
        ram_cell[    2244] = 32'h00000000;
        ram_cell[    2245] = 32'h00000000;
        ram_cell[    2246] = 32'h00000000;
        ram_cell[    2247] = 32'h00000000;
        ram_cell[    2248] = 32'h00000000;
        ram_cell[    2249] = 32'h00000000;
        ram_cell[    2250] = 32'h00000000;
        ram_cell[    2251] = 32'h00000000;
        ram_cell[    2252] = 32'h00000000;
        ram_cell[    2253] = 32'h00000000;
        ram_cell[    2254] = 32'h00000000;
        ram_cell[    2255] = 32'h00000000;
        ram_cell[    2256] = 32'h00000000;
        ram_cell[    2257] = 32'h00000000;
        ram_cell[    2258] = 32'h00000000;
        ram_cell[    2259] = 32'h00000000;
        ram_cell[    2260] = 32'h00000000;
        ram_cell[    2261] = 32'h00000000;
        ram_cell[    2262] = 32'h00000000;
        ram_cell[    2263] = 32'h00000000;
        ram_cell[    2264] = 32'h00000000;
        ram_cell[    2265] = 32'h00000000;
        ram_cell[    2266] = 32'h00000000;
        ram_cell[    2267] = 32'h00000000;
        ram_cell[    2268] = 32'h00000000;
        ram_cell[    2269] = 32'h00000000;
        ram_cell[    2270] = 32'h00000000;
        ram_cell[    2271] = 32'h00000000;
        ram_cell[    2272] = 32'h00000000;
        ram_cell[    2273] = 32'h00000000;
        ram_cell[    2274] = 32'h00000000;
        ram_cell[    2275] = 32'h00000000;
        ram_cell[    2276] = 32'h00000000;
        ram_cell[    2277] = 32'h00000000;
        ram_cell[    2278] = 32'h00000000;
        ram_cell[    2279] = 32'h00000000;
        ram_cell[    2280] = 32'h00000000;
        ram_cell[    2281] = 32'h00000000;
        ram_cell[    2282] = 32'h00000000;
        ram_cell[    2283] = 32'h00000000;
        ram_cell[    2284] = 32'h00000000;
        ram_cell[    2285] = 32'h00000000;
        ram_cell[    2286] = 32'h00000000;
        ram_cell[    2287] = 32'h00000000;
        ram_cell[    2288] = 32'h00000000;
        ram_cell[    2289] = 32'h00000000;
        ram_cell[    2290] = 32'h00000000;
        ram_cell[    2291] = 32'h00000000;
        ram_cell[    2292] = 32'h00000000;
        ram_cell[    2293] = 32'h00000000;
        ram_cell[    2294] = 32'h00000000;
        ram_cell[    2295] = 32'h00000000;
        ram_cell[    2296] = 32'h00000000;
        ram_cell[    2297] = 32'h00000000;
        ram_cell[    2298] = 32'h00000000;
        ram_cell[    2299] = 32'h00000000;
        ram_cell[    2300] = 32'h00000000;
        ram_cell[    2301] = 32'h00000000;
        ram_cell[    2302] = 32'h00000000;
        ram_cell[    2303] = 32'h00000000;
        ram_cell[    2304] = 32'h00000000;
        ram_cell[    2305] = 32'h00000000;
        ram_cell[    2306] = 32'h00000000;
        ram_cell[    2307] = 32'h00000000;
        ram_cell[    2308] = 32'h00000000;
        ram_cell[    2309] = 32'h00000000;
        ram_cell[    2310] = 32'h00000000;
        ram_cell[    2311] = 32'h00000000;
        ram_cell[    2312] = 32'h00000000;
        ram_cell[    2313] = 32'h00000000;
        ram_cell[    2314] = 32'h00000000;
        ram_cell[    2315] = 32'h00000000;
        ram_cell[    2316] = 32'h00000000;
        ram_cell[    2317] = 32'h00000000;
        ram_cell[    2318] = 32'h00000000;
        ram_cell[    2319] = 32'h00000000;
        ram_cell[    2320] = 32'h00000000;
        ram_cell[    2321] = 32'h00000000;
        ram_cell[    2322] = 32'h00000000;
        ram_cell[    2323] = 32'h00000000;
        ram_cell[    2324] = 32'h00000000;
        ram_cell[    2325] = 32'h00000000;
        ram_cell[    2326] = 32'h00000000;
        ram_cell[    2327] = 32'h00000000;
        ram_cell[    2328] = 32'h00000000;
        ram_cell[    2329] = 32'h00000000;
        ram_cell[    2330] = 32'h00000000;
        ram_cell[    2331] = 32'h00000000;
        ram_cell[    2332] = 32'h00000000;
        ram_cell[    2333] = 32'h00000000;
        ram_cell[    2334] = 32'h00000000;
        ram_cell[    2335] = 32'h00000000;
        ram_cell[    2336] = 32'h00000000;
        ram_cell[    2337] = 32'h00000000;
        ram_cell[    2338] = 32'h00000000;
        ram_cell[    2339] = 32'h00000000;
        ram_cell[    2340] = 32'h00000000;
        ram_cell[    2341] = 32'h00000000;
        ram_cell[    2342] = 32'h00000000;
        ram_cell[    2343] = 32'h00000000;
        ram_cell[    2344] = 32'h00000000;
        ram_cell[    2345] = 32'h00000000;
        ram_cell[    2346] = 32'h00000000;
        ram_cell[    2347] = 32'h00000000;
        ram_cell[    2348] = 32'h00000000;
        ram_cell[    2349] = 32'h00000000;
        ram_cell[    2350] = 32'h00000000;
        ram_cell[    2351] = 32'h00000000;
        ram_cell[    2352] = 32'h00000000;
        ram_cell[    2353] = 32'h00000000;
        ram_cell[    2354] = 32'h00000000;
        ram_cell[    2355] = 32'h00000000;
        ram_cell[    2356] = 32'h00000000;
        ram_cell[    2357] = 32'h00000000;
        ram_cell[    2358] = 32'h00000000;
        ram_cell[    2359] = 32'h00000000;
        ram_cell[    2360] = 32'h00000000;
        ram_cell[    2361] = 32'h00000000;
        ram_cell[    2362] = 32'h00000000;
        ram_cell[    2363] = 32'h00000000;
        ram_cell[    2364] = 32'h00000000;
        ram_cell[    2365] = 32'h00000000;
        ram_cell[    2366] = 32'h00000000;
        ram_cell[    2367] = 32'h00000000;
        ram_cell[    2368] = 32'h00000000;
        ram_cell[    2369] = 32'h00000000;
        ram_cell[    2370] = 32'h00000000;
        ram_cell[    2371] = 32'h00000000;
        ram_cell[    2372] = 32'h00000000;
        ram_cell[    2373] = 32'h00000000;
        ram_cell[    2374] = 32'h00000000;
        ram_cell[    2375] = 32'h00000000;
        ram_cell[    2376] = 32'h00000000;
        ram_cell[    2377] = 32'h00000000;
        ram_cell[    2378] = 32'h00000000;
        ram_cell[    2379] = 32'h00000000;
        ram_cell[    2380] = 32'h00000000;
        ram_cell[    2381] = 32'h00000000;
        ram_cell[    2382] = 32'h00000000;
        ram_cell[    2383] = 32'h00000000;
        ram_cell[    2384] = 32'h00000000;
        ram_cell[    2385] = 32'h00000000;
        ram_cell[    2386] = 32'h00000000;
        ram_cell[    2387] = 32'h00000000;
        ram_cell[    2388] = 32'h00000000;
        ram_cell[    2389] = 32'h00000000;
        ram_cell[    2390] = 32'h00000000;
        ram_cell[    2391] = 32'h00000000;
        ram_cell[    2392] = 32'h00000000;
        ram_cell[    2393] = 32'h00000000;
        ram_cell[    2394] = 32'h00000000;
        ram_cell[    2395] = 32'h00000000;
        ram_cell[    2396] = 32'h00000000;
        ram_cell[    2397] = 32'h00000000;
        ram_cell[    2398] = 32'h00000000;
        ram_cell[    2399] = 32'h00000000;
        ram_cell[    2400] = 32'h00000000;
        ram_cell[    2401] = 32'h00000000;
        ram_cell[    2402] = 32'h00000000;
        ram_cell[    2403] = 32'h00000000;
        ram_cell[    2404] = 32'h00000000;
        ram_cell[    2405] = 32'h00000000;
        ram_cell[    2406] = 32'h00000000;
        ram_cell[    2407] = 32'h00000000;
        ram_cell[    2408] = 32'h00000000;
        ram_cell[    2409] = 32'h00000000;
        ram_cell[    2410] = 32'h00000000;
        ram_cell[    2411] = 32'h00000000;
        ram_cell[    2412] = 32'h00000000;
        ram_cell[    2413] = 32'h00000000;
        ram_cell[    2414] = 32'h00000000;
        ram_cell[    2415] = 32'h00000000;
        ram_cell[    2416] = 32'h00000000;
        ram_cell[    2417] = 32'h00000000;
        ram_cell[    2418] = 32'h00000000;
        ram_cell[    2419] = 32'h00000000;
        ram_cell[    2420] = 32'h00000000;
        ram_cell[    2421] = 32'h00000000;
        ram_cell[    2422] = 32'h00000000;
        ram_cell[    2423] = 32'h00000000;
        ram_cell[    2424] = 32'h00000000;
        ram_cell[    2425] = 32'h00000000;
        ram_cell[    2426] = 32'h00000000;
        ram_cell[    2427] = 32'h00000000;
        ram_cell[    2428] = 32'h00000000;
        ram_cell[    2429] = 32'h00000000;
        ram_cell[    2430] = 32'h00000000;
        ram_cell[    2431] = 32'h00000000;
        ram_cell[    2432] = 32'h00000000;
        ram_cell[    2433] = 32'h00000000;
        ram_cell[    2434] = 32'h00000000;
        ram_cell[    2435] = 32'h00000000;
        ram_cell[    2436] = 32'h00000000;
        ram_cell[    2437] = 32'h00000000;
        ram_cell[    2438] = 32'h00000000;
        ram_cell[    2439] = 32'h00000000;
        ram_cell[    2440] = 32'h00000000;
        ram_cell[    2441] = 32'h00000000;
        ram_cell[    2442] = 32'h00000000;
        ram_cell[    2443] = 32'h00000000;
        ram_cell[    2444] = 32'h00000000;
        ram_cell[    2445] = 32'h00000000;
        ram_cell[    2446] = 32'h00000000;
        ram_cell[    2447] = 32'h00000000;
        ram_cell[    2448] = 32'h00000000;
        ram_cell[    2449] = 32'h00000000;
        ram_cell[    2450] = 32'h00000000;
        ram_cell[    2451] = 32'h00000000;
        ram_cell[    2452] = 32'h00000000;
        ram_cell[    2453] = 32'h00000000;
        ram_cell[    2454] = 32'h00000000;
        ram_cell[    2455] = 32'h00000000;
        ram_cell[    2456] = 32'h00000000;
        ram_cell[    2457] = 32'h00000000;
        ram_cell[    2458] = 32'h00000000;
        ram_cell[    2459] = 32'h00000000;
        ram_cell[    2460] = 32'h00000000;
        ram_cell[    2461] = 32'h00000000;
        ram_cell[    2462] = 32'h00000000;
        ram_cell[    2463] = 32'h00000000;
        ram_cell[    2464] = 32'h00000000;
        ram_cell[    2465] = 32'h00000000;
        ram_cell[    2466] = 32'h00000000;
        ram_cell[    2467] = 32'h00000000;
        ram_cell[    2468] = 32'h00000000;
        ram_cell[    2469] = 32'h00000000;
        ram_cell[    2470] = 32'h00000000;
        ram_cell[    2471] = 32'h00000000;
        ram_cell[    2472] = 32'h00000000;
        ram_cell[    2473] = 32'h00000000;
        ram_cell[    2474] = 32'h00000000;
        ram_cell[    2475] = 32'h00000000;
        ram_cell[    2476] = 32'h00000000;
        ram_cell[    2477] = 32'h00000000;
        ram_cell[    2478] = 32'h00000000;
        ram_cell[    2479] = 32'h00000000;
        ram_cell[    2480] = 32'h00000000;
        ram_cell[    2481] = 32'h00000000;
        ram_cell[    2482] = 32'h00000000;
        ram_cell[    2483] = 32'h00000000;
        ram_cell[    2484] = 32'h00000000;
        ram_cell[    2485] = 32'h00000000;
        ram_cell[    2486] = 32'h00000000;
        ram_cell[    2487] = 32'h00000000;
        ram_cell[    2488] = 32'h00000000;
        ram_cell[    2489] = 32'h00000000;
        ram_cell[    2490] = 32'h00000000;
        ram_cell[    2491] = 32'h00000000;
        ram_cell[    2492] = 32'h00000000;
        ram_cell[    2493] = 32'h00000000;
        ram_cell[    2494] = 32'h00000000;
        ram_cell[    2495] = 32'h00000000;
        ram_cell[    2496] = 32'h00000000;
        ram_cell[    2497] = 32'h00000000;
        ram_cell[    2498] = 32'h00000000;
        ram_cell[    2499] = 32'h00000000;
        ram_cell[    2500] = 32'h00000000;
        ram_cell[    2501] = 32'h00000000;
        ram_cell[    2502] = 32'h00000000;
        ram_cell[    2503] = 32'h00000000;
        ram_cell[    2504] = 32'h00000000;
        ram_cell[    2505] = 32'h00000000;
        ram_cell[    2506] = 32'h00000000;
        ram_cell[    2507] = 32'h00000000;
        ram_cell[    2508] = 32'h00000000;
        ram_cell[    2509] = 32'h00000000;
        ram_cell[    2510] = 32'h00000000;
        ram_cell[    2511] = 32'h00000000;
        ram_cell[    2512] = 32'h00000000;
        ram_cell[    2513] = 32'h00000000;
        ram_cell[    2514] = 32'h00000000;
        ram_cell[    2515] = 32'h00000000;
        ram_cell[    2516] = 32'h00000000;
        ram_cell[    2517] = 32'h00000000;
        ram_cell[    2518] = 32'h00000000;
        ram_cell[    2519] = 32'h00000000;
        ram_cell[    2520] = 32'h00000000;
        ram_cell[    2521] = 32'h00000000;
        ram_cell[    2522] = 32'h00000000;
        ram_cell[    2523] = 32'h00000000;
        ram_cell[    2524] = 32'h00000000;
        ram_cell[    2525] = 32'h00000000;
        ram_cell[    2526] = 32'h00000000;
        ram_cell[    2527] = 32'h00000000;
        ram_cell[    2528] = 32'h00000000;
        ram_cell[    2529] = 32'h00000000;
        ram_cell[    2530] = 32'h00000000;
        ram_cell[    2531] = 32'h00000000;
        ram_cell[    2532] = 32'h00000000;
        ram_cell[    2533] = 32'h00000000;
        ram_cell[    2534] = 32'h00000000;
        ram_cell[    2535] = 32'h00000000;
        ram_cell[    2536] = 32'h00000000;
        ram_cell[    2537] = 32'h00000000;
        ram_cell[    2538] = 32'h00000000;
        ram_cell[    2539] = 32'h00000000;
        ram_cell[    2540] = 32'h00000000;
        ram_cell[    2541] = 32'h00000000;
        ram_cell[    2542] = 32'h00000000;
        ram_cell[    2543] = 32'h00000000;
        ram_cell[    2544] = 32'h00000000;
        ram_cell[    2545] = 32'h00000000;
        ram_cell[    2546] = 32'h00000000;
        ram_cell[    2547] = 32'h00000000;
        ram_cell[    2548] = 32'h00000000;
        ram_cell[    2549] = 32'h00000000;
        ram_cell[    2550] = 32'h00000000;
        ram_cell[    2551] = 32'h00000000;
        ram_cell[    2552] = 32'h00000000;
        ram_cell[    2553] = 32'h00000000;
        ram_cell[    2554] = 32'h00000000;
        ram_cell[    2555] = 32'h00000000;
        ram_cell[    2556] = 32'h00000000;
        ram_cell[    2557] = 32'h00000000;
        ram_cell[    2558] = 32'h00000000;
        ram_cell[    2559] = 32'h00000000;
        ram_cell[    2560] = 32'h00000000;
        ram_cell[    2561] = 32'h00000000;
        ram_cell[    2562] = 32'h00000000;
        ram_cell[    2563] = 32'h00000000;
        ram_cell[    2564] = 32'h00000000;
        ram_cell[    2565] = 32'h00000000;
        ram_cell[    2566] = 32'h00000000;
        ram_cell[    2567] = 32'h00000000;
        ram_cell[    2568] = 32'h00000000;
        ram_cell[    2569] = 32'h00000000;
        ram_cell[    2570] = 32'h00000000;
        ram_cell[    2571] = 32'h00000000;
        ram_cell[    2572] = 32'h00000000;
        ram_cell[    2573] = 32'h00000000;
        ram_cell[    2574] = 32'h00000000;
        ram_cell[    2575] = 32'h00000000;
        ram_cell[    2576] = 32'h00000000;
        ram_cell[    2577] = 32'h00000000;
        ram_cell[    2578] = 32'h00000000;
        ram_cell[    2579] = 32'h00000000;
        ram_cell[    2580] = 32'h00000000;
        ram_cell[    2581] = 32'h00000000;
        ram_cell[    2582] = 32'h00000000;
        ram_cell[    2583] = 32'h00000000;
        ram_cell[    2584] = 32'h00000000;
        ram_cell[    2585] = 32'h00000000;
        ram_cell[    2586] = 32'h00000000;
        ram_cell[    2587] = 32'h00000000;
        ram_cell[    2588] = 32'h00000000;
        ram_cell[    2589] = 32'h00000000;
        ram_cell[    2590] = 32'h00000000;
        ram_cell[    2591] = 32'h00000000;
        ram_cell[    2592] = 32'h00000000;
        ram_cell[    2593] = 32'h00000000;
        ram_cell[    2594] = 32'h00000000;
        ram_cell[    2595] = 32'h00000000;
        ram_cell[    2596] = 32'h00000000;
        ram_cell[    2597] = 32'h00000000;
        ram_cell[    2598] = 32'h00000000;
        ram_cell[    2599] = 32'h00000000;
        ram_cell[    2600] = 32'h00000000;
        ram_cell[    2601] = 32'h00000000;
        ram_cell[    2602] = 32'h00000000;
        ram_cell[    2603] = 32'h00000000;
        ram_cell[    2604] = 32'h00000000;
        ram_cell[    2605] = 32'h00000000;
        ram_cell[    2606] = 32'h00000000;
        ram_cell[    2607] = 32'h00000000;
        ram_cell[    2608] = 32'h00000000;
        ram_cell[    2609] = 32'h00000000;
        ram_cell[    2610] = 32'h00000000;
        ram_cell[    2611] = 32'h00000000;
        ram_cell[    2612] = 32'h00000000;
        ram_cell[    2613] = 32'h00000000;
        ram_cell[    2614] = 32'h00000000;
        ram_cell[    2615] = 32'h00000000;
        ram_cell[    2616] = 32'h00000000;
        ram_cell[    2617] = 32'h00000000;
        ram_cell[    2618] = 32'h00000000;
        ram_cell[    2619] = 32'h00000000;
        ram_cell[    2620] = 32'h00000000;
        ram_cell[    2621] = 32'h00000000;
        ram_cell[    2622] = 32'h00000000;
        ram_cell[    2623] = 32'h00000000;
        ram_cell[    2624] = 32'h00000000;
        ram_cell[    2625] = 32'h00000000;
        ram_cell[    2626] = 32'h00000000;
        ram_cell[    2627] = 32'h00000000;
        ram_cell[    2628] = 32'h00000000;
        ram_cell[    2629] = 32'h00000000;
        ram_cell[    2630] = 32'h00000000;
        ram_cell[    2631] = 32'h00000000;
        ram_cell[    2632] = 32'h00000000;
        ram_cell[    2633] = 32'h00000000;
        ram_cell[    2634] = 32'h00000000;
        ram_cell[    2635] = 32'h00000000;
        ram_cell[    2636] = 32'h00000000;
        ram_cell[    2637] = 32'h00000000;
        ram_cell[    2638] = 32'h00000000;
        ram_cell[    2639] = 32'h00000000;
        ram_cell[    2640] = 32'h00000000;
        ram_cell[    2641] = 32'h00000000;
        ram_cell[    2642] = 32'h00000000;
        ram_cell[    2643] = 32'h00000000;
        ram_cell[    2644] = 32'h00000000;
        ram_cell[    2645] = 32'h00000000;
        ram_cell[    2646] = 32'h00000000;
        ram_cell[    2647] = 32'h00000000;
        ram_cell[    2648] = 32'h00000000;
        ram_cell[    2649] = 32'h00000000;
        ram_cell[    2650] = 32'h00000000;
        ram_cell[    2651] = 32'h00000000;
        ram_cell[    2652] = 32'h00000000;
        ram_cell[    2653] = 32'h00000000;
        ram_cell[    2654] = 32'h00000000;
        ram_cell[    2655] = 32'h00000000;
        ram_cell[    2656] = 32'h00000000;
        ram_cell[    2657] = 32'h00000000;
        ram_cell[    2658] = 32'h00000000;
        ram_cell[    2659] = 32'h00000000;
        ram_cell[    2660] = 32'h00000000;
        ram_cell[    2661] = 32'h00000000;
        ram_cell[    2662] = 32'h00000000;
        ram_cell[    2663] = 32'h00000000;
        ram_cell[    2664] = 32'h00000000;
        ram_cell[    2665] = 32'h00000000;
        ram_cell[    2666] = 32'h00000000;
        ram_cell[    2667] = 32'h00000000;
        ram_cell[    2668] = 32'h00000000;
        ram_cell[    2669] = 32'h00000000;
        ram_cell[    2670] = 32'h00000000;
        ram_cell[    2671] = 32'h00000000;
        ram_cell[    2672] = 32'h00000000;
        ram_cell[    2673] = 32'h00000000;
        ram_cell[    2674] = 32'h00000000;
        ram_cell[    2675] = 32'h00000000;
        ram_cell[    2676] = 32'h00000000;
        ram_cell[    2677] = 32'h00000000;
        ram_cell[    2678] = 32'h00000000;
        ram_cell[    2679] = 32'h00000000;
        ram_cell[    2680] = 32'h00000000;
        ram_cell[    2681] = 32'h00000000;
        ram_cell[    2682] = 32'h00000000;
        ram_cell[    2683] = 32'h00000000;
        ram_cell[    2684] = 32'h00000000;
        ram_cell[    2685] = 32'h00000000;
        ram_cell[    2686] = 32'h00000000;
        ram_cell[    2687] = 32'h00000000;
        ram_cell[    2688] = 32'h00000000;
        ram_cell[    2689] = 32'h00000000;
        ram_cell[    2690] = 32'h00000000;
        ram_cell[    2691] = 32'h00000000;
        ram_cell[    2692] = 32'h00000000;
        ram_cell[    2693] = 32'h00000000;
        ram_cell[    2694] = 32'h00000000;
        ram_cell[    2695] = 32'h00000000;
        ram_cell[    2696] = 32'h00000000;
        ram_cell[    2697] = 32'h00000000;
        ram_cell[    2698] = 32'h00000000;
        ram_cell[    2699] = 32'h00000000;
        ram_cell[    2700] = 32'h00000000;
        ram_cell[    2701] = 32'h00000000;
        ram_cell[    2702] = 32'h00000000;
        ram_cell[    2703] = 32'h00000000;
        ram_cell[    2704] = 32'h00000000;
        ram_cell[    2705] = 32'h00000000;
        ram_cell[    2706] = 32'h00000000;
        ram_cell[    2707] = 32'h00000000;
        ram_cell[    2708] = 32'h00000000;
        ram_cell[    2709] = 32'h00000000;
        ram_cell[    2710] = 32'h00000000;
        ram_cell[    2711] = 32'h00000000;
        ram_cell[    2712] = 32'h00000000;
        ram_cell[    2713] = 32'h00000000;
        ram_cell[    2714] = 32'h00000000;
        ram_cell[    2715] = 32'h00000000;
        ram_cell[    2716] = 32'h00000000;
        ram_cell[    2717] = 32'h00000000;
        ram_cell[    2718] = 32'h00000000;
        ram_cell[    2719] = 32'h00000000;
        ram_cell[    2720] = 32'h00000000;
        ram_cell[    2721] = 32'h00000000;
        ram_cell[    2722] = 32'h00000000;
        ram_cell[    2723] = 32'h00000000;
        ram_cell[    2724] = 32'h00000000;
        ram_cell[    2725] = 32'h00000000;
        ram_cell[    2726] = 32'h00000000;
        ram_cell[    2727] = 32'h00000000;
        ram_cell[    2728] = 32'h00000000;
        ram_cell[    2729] = 32'h00000000;
        ram_cell[    2730] = 32'h00000000;
        ram_cell[    2731] = 32'h00000000;
        ram_cell[    2732] = 32'h00000000;
        ram_cell[    2733] = 32'h00000000;
        ram_cell[    2734] = 32'h00000000;
        ram_cell[    2735] = 32'h00000000;
        ram_cell[    2736] = 32'h00000000;
        ram_cell[    2737] = 32'h00000000;
        ram_cell[    2738] = 32'h00000000;
        ram_cell[    2739] = 32'h00000000;
        ram_cell[    2740] = 32'h00000000;
        ram_cell[    2741] = 32'h00000000;
        ram_cell[    2742] = 32'h00000000;
        ram_cell[    2743] = 32'h00000000;
        ram_cell[    2744] = 32'h00000000;
        ram_cell[    2745] = 32'h00000000;
        ram_cell[    2746] = 32'h00000000;
        ram_cell[    2747] = 32'h00000000;
        ram_cell[    2748] = 32'h00000000;
        ram_cell[    2749] = 32'h00000000;
        ram_cell[    2750] = 32'h00000000;
        ram_cell[    2751] = 32'h00000000;
        ram_cell[    2752] = 32'h00000000;
        ram_cell[    2753] = 32'h00000000;
        ram_cell[    2754] = 32'h00000000;
        ram_cell[    2755] = 32'h00000000;
        ram_cell[    2756] = 32'h00000000;
        ram_cell[    2757] = 32'h00000000;
        ram_cell[    2758] = 32'h00000000;
        ram_cell[    2759] = 32'h00000000;
        ram_cell[    2760] = 32'h00000000;
        ram_cell[    2761] = 32'h00000000;
        ram_cell[    2762] = 32'h00000000;
        ram_cell[    2763] = 32'h00000000;
        ram_cell[    2764] = 32'h00000000;
        ram_cell[    2765] = 32'h00000000;
        ram_cell[    2766] = 32'h00000000;
        ram_cell[    2767] = 32'h00000000;
        ram_cell[    2768] = 32'h00000000;
        ram_cell[    2769] = 32'h00000000;
        ram_cell[    2770] = 32'h00000000;
        ram_cell[    2771] = 32'h00000000;
        ram_cell[    2772] = 32'h00000000;
        ram_cell[    2773] = 32'h00000000;
        ram_cell[    2774] = 32'h00000000;
        ram_cell[    2775] = 32'h00000000;
        ram_cell[    2776] = 32'h00000000;
        ram_cell[    2777] = 32'h00000000;
        ram_cell[    2778] = 32'h00000000;
        ram_cell[    2779] = 32'h00000000;
        ram_cell[    2780] = 32'h00000000;
        ram_cell[    2781] = 32'h00000000;
        ram_cell[    2782] = 32'h00000000;
        ram_cell[    2783] = 32'h00000000;
        ram_cell[    2784] = 32'h00000000;
        ram_cell[    2785] = 32'h00000000;
        ram_cell[    2786] = 32'h00000000;
        ram_cell[    2787] = 32'h00000000;
        ram_cell[    2788] = 32'h00000000;
        ram_cell[    2789] = 32'h00000000;
        ram_cell[    2790] = 32'h00000000;
        ram_cell[    2791] = 32'h00000000;
        ram_cell[    2792] = 32'h00000000;
        ram_cell[    2793] = 32'h00000000;
        ram_cell[    2794] = 32'h00000000;
        ram_cell[    2795] = 32'h00000000;
        ram_cell[    2796] = 32'h00000000;
        ram_cell[    2797] = 32'h00000000;
        ram_cell[    2798] = 32'h00000000;
        ram_cell[    2799] = 32'h00000000;
        ram_cell[    2800] = 32'h00000000;
        ram_cell[    2801] = 32'h00000000;
        ram_cell[    2802] = 32'h00000000;
        ram_cell[    2803] = 32'h00000000;
        ram_cell[    2804] = 32'h00000000;
        ram_cell[    2805] = 32'h00000000;
        ram_cell[    2806] = 32'h00000000;
        ram_cell[    2807] = 32'h00000000;
        ram_cell[    2808] = 32'h00000000;
        ram_cell[    2809] = 32'h00000000;
        ram_cell[    2810] = 32'h00000000;
        ram_cell[    2811] = 32'h00000000;
        ram_cell[    2812] = 32'h00000000;
        ram_cell[    2813] = 32'h00000000;
        ram_cell[    2814] = 32'h00000000;
        ram_cell[    2815] = 32'h00000000;
        ram_cell[    2816] = 32'h00000000;
        ram_cell[    2817] = 32'h00000000;
        ram_cell[    2818] = 32'h00000000;
        ram_cell[    2819] = 32'h00000000;
        ram_cell[    2820] = 32'h00000000;
        ram_cell[    2821] = 32'h00000000;
        ram_cell[    2822] = 32'h00000000;
        ram_cell[    2823] = 32'h00000000;
        ram_cell[    2824] = 32'h00000000;
        ram_cell[    2825] = 32'h00000000;
        ram_cell[    2826] = 32'h00000000;
        ram_cell[    2827] = 32'h00000000;
        ram_cell[    2828] = 32'h00000000;
        ram_cell[    2829] = 32'h00000000;
        ram_cell[    2830] = 32'h00000000;
        ram_cell[    2831] = 32'h00000000;
        ram_cell[    2832] = 32'h00000000;
        ram_cell[    2833] = 32'h00000000;
        ram_cell[    2834] = 32'h00000000;
        ram_cell[    2835] = 32'h00000000;
        ram_cell[    2836] = 32'h00000000;
        ram_cell[    2837] = 32'h00000000;
        ram_cell[    2838] = 32'h00000000;
        ram_cell[    2839] = 32'h00000000;
        ram_cell[    2840] = 32'h00000000;
        ram_cell[    2841] = 32'h00000000;
        ram_cell[    2842] = 32'h00000000;
        ram_cell[    2843] = 32'h00000000;
        ram_cell[    2844] = 32'h00000000;
        ram_cell[    2845] = 32'h00000000;
        ram_cell[    2846] = 32'h00000000;
        ram_cell[    2847] = 32'h00000000;
        ram_cell[    2848] = 32'h00000000;
        ram_cell[    2849] = 32'h00000000;
        ram_cell[    2850] = 32'h00000000;
        ram_cell[    2851] = 32'h00000000;
        ram_cell[    2852] = 32'h00000000;
        ram_cell[    2853] = 32'h00000000;
        ram_cell[    2854] = 32'h00000000;
        ram_cell[    2855] = 32'h00000000;
        ram_cell[    2856] = 32'h00000000;
        ram_cell[    2857] = 32'h00000000;
        ram_cell[    2858] = 32'h00000000;
        ram_cell[    2859] = 32'h00000000;
        ram_cell[    2860] = 32'h00000000;
        ram_cell[    2861] = 32'h00000000;
        ram_cell[    2862] = 32'h00000000;
        ram_cell[    2863] = 32'h00000000;
        ram_cell[    2864] = 32'h00000000;
        ram_cell[    2865] = 32'h00000000;
        ram_cell[    2866] = 32'h00000000;
        ram_cell[    2867] = 32'h00000000;
        ram_cell[    2868] = 32'h00000000;
        ram_cell[    2869] = 32'h00000000;
        ram_cell[    2870] = 32'h00000000;
        ram_cell[    2871] = 32'h00000000;
        ram_cell[    2872] = 32'h00000000;
        ram_cell[    2873] = 32'h00000000;
        ram_cell[    2874] = 32'h00000000;
        ram_cell[    2875] = 32'h00000000;
        ram_cell[    2876] = 32'h00000000;
        ram_cell[    2877] = 32'h00000000;
        ram_cell[    2878] = 32'h00000000;
        ram_cell[    2879] = 32'h00000000;
        ram_cell[    2880] = 32'h00000000;
        ram_cell[    2881] = 32'h00000000;
        ram_cell[    2882] = 32'h00000000;
        ram_cell[    2883] = 32'h00000000;
        ram_cell[    2884] = 32'h00000000;
        ram_cell[    2885] = 32'h00000000;
        ram_cell[    2886] = 32'h00000000;
        ram_cell[    2887] = 32'h00000000;
        ram_cell[    2888] = 32'h00000000;
        ram_cell[    2889] = 32'h00000000;
        ram_cell[    2890] = 32'h00000000;
        ram_cell[    2891] = 32'h00000000;
        ram_cell[    2892] = 32'h00000000;
        ram_cell[    2893] = 32'h00000000;
        ram_cell[    2894] = 32'h00000000;
        ram_cell[    2895] = 32'h00000000;
        ram_cell[    2896] = 32'h00000000;
        ram_cell[    2897] = 32'h00000000;
        ram_cell[    2898] = 32'h00000000;
        ram_cell[    2899] = 32'h00000000;
        ram_cell[    2900] = 32'h00000000;
        ram_cell[    2901] = 32'h00000000;
        ram_cell[    2902] = 32'h00000000;
        ram_cell[    2903] = 32'h00000000;
        ram_cell[    2904] = 32'h00000000;
        ram_cell[    2905] = 32'h00000000;
        ram_cell[    2906] = 32'h00000000;
        ram_cell[    2907] = 32'h00000000;
        ram_cell[    2908] = 32'h00000000;
        ram_cell[    2909] = 32'h00000000;
        ram_cell[    2910] = 32'h00000000;
        ram_cell[    2911] = 32'h00000000;
        ram_cell[    2912] = 32'h00000000;
        ram_cell[    2913] = 32'h00000000;
        ram_cell[    2914] = 32'h00000000;
        ram_cell[    2915] = 32'h00000000;
        ram_cell[    2916] = 32'h00000000;
        ram_cell[    2917] = 32'h00000000;
        ram_cell[    2918] = 32'h00000000;
        ram_cell[    2919] = 32'h00000000;
        ram_cell[    2920] = 32'h00000000;
        ram_cell[    2921] = 32'h00000000;
        ram_cell[    2922] = 32'h00000000;
        ram_cell[    2923] = 32'h00000000;
        ram_cell[    2924] = 32'h00000000;
        ram_cell[    2925] = 32'h00000000;
        ram_cell[    2926] = 32'h00000000;
        ram_cell[    2927] = 32'h00000000;
        ram_cell[    2928] = 32'h00000000;
        ram_cell[    2929] = 32'h00000000;
        ram_cell[    2930] = 32'h00000000;
        ram_cell[    2931] = 32'h00000000;
        ram_cell[    2932] = 32'h00000000;
        ram_cell[    2933] = 32'h00000000;
        ram_cell[    2934] = 32'h00000000;
        ram_cell[    2935] = 32'h00000000;
        ram_cell[    2936] = 32'h00000000;
        ram_cell[    2937] = 32'h00000000;
        ram_cell[    2938] = 32'h00000000;
        ram_cell[    2939] = 32'h00000000;
        ram_cell[    2940] = 32'h00000000;
        ram_cell[    2941] = 32'h00000000;
        ram_cell[    2942] = 32'h00000000;
        ram_cell[    2943] = 32'h00000000;
        ram_cell[    2944] = 32'h00000000;
        ram_cell[    2945] = 32'h00000000;
        ram_cell[    2946] = 32'h00000000;
        ram_cell[    2947] = 32'h00000000;
        ram_cell[    2948] = 32'h00000000;
        ram_cell[    2949] = 32'h00000000;
        ram_cell[    2950] = 32'h00000000;
        ram_cell[    2951] = 32'h00000000;
        ram_cell[    2952] = 32'h00000000;
        ram_cell[    2953] = 32'h00000000;
        ram_cell[    2954] = 32'h00000000;
        ram_cell[    2955] = 32'h00000000;
        ram_cell[    2956] = 32'h00000000;
        ram_cell[    2957] = 32'h00000000;
        ram_cell[    2958] = 32'h00000000;
        ram_cell[    2959] = 32'h00000000;
        ram_cell[    2960] = 32'h00000000;
        ram_cell[    2961] = 32'h00000000;
        ram_cell[    2962] = 32'h00000000;
        ram_cell[    2963] = 32'h00000000;
        ram_cell[    2964] = 32'h00000000;
        ram_cell[    2965] = 32'h00000000;
        ram_cell[    2966] = 32'h00000000;
        ram_cell[    2967] = 32'h00000000;
        ram_cell[    2968] = 32'h00000000;
        ram_cell[    2969] = 32'h00000000;
        ram_cell[    2970] = 32'h00000000;
        ram_cell[    2971] = 32'h00000000;
        ram_cell[    2972] = 32'h00000000;
        ram_cell[    2973] = 32'h00000000;
        ram_cell[    2974] = 32'h00000000;
        ram_cell[    2975] = 32'h00000000;
        ram_cell[    2976] = 32'h00000000;
        ram_cell[    2977] = 32'h00000000;
        ram_cell[    2978] = 32'h00000000;
        ram_cell[    2979] = 32'h00000000;
        ram_cell[    2980] = 32'h00000000;
        ram_cell[    2981] = 32'h00000000;
        ram_cell[    2982] = 32'h00000000;
        ram_cell[    2983] = 32'h00000000;
        ram_cell[    2984] = 32'h00000000;
        ram_cell[    2985] = 32'h00000000;
        ram_cell[    2986] = 32'h00000000;
        ram_cell[    2987] = 32'h00000000;
        ram_cell[    2988] = 32'h00000000;
        ram_cell[    2989] = 32'h00000000;
        ram_cell[    2990] = 32'h00000000;
        ram_cell[    2991] = 32'h00000000;
        ram_cell[    2992] = 32'h00000000;
        ram_cell[    2993] = 32'h00000000;
        ram_cell[    2994] = 32'h00000000;
        ram_cell[    2995] = 32'h00000000;
        ram_cell[    2996] = 32'h00000000;
        ram_cell[    2997] = 32'h00000000;
        ram_cell[    2998] = 32'h00000000;
        ram_cell[    2999] = 32'h00000000;
        ram_cell[    3000] = 32'h00000000;
        ram_cell[    3001] = 32'h00000000;
        ram_cell[    3002] = 32'h00000000;
        ram_cell[    3003] = 32'h00000000;
        ram_cell[    3004] = 32'h00000000;
        ram_cell[    3005] = 32'h00000000;
        ram_cell[    3006] = 32'h00000000;
        ram_cell[    3007] = 32'h00000000;
        ram_cell[    3008] = 32'h00000000;
        ram_cell[    3009] = 32'h00000000;
        ram_cell[    3010] = 32'h00000000;
        ram_cell[    3011] = 32'h00000000;
        ram_cell[    3012] = 32'h00000000;
        ram_cell[    3013] = 32'h00000000;
        ram_cell[    3014] = 32'h00000000;
        ram_cell[    3015] = 32'h00000000;
        ram_cell[    3016] = 32'h00000000;
        ram_cell[    3017] = 32'h00000000;
        ram_cell[    3018] = 32'h00000000;
        ram_cell[    3019] = 32'h00000000;
        ram_cell[    3020] = 32'h00000000;
        ram_cell[    3021] = 32'h00000000;
        ram_cell[    3022] = 32'h00000000;
        ram_cell[    3023] = 32'h00000000;
        ram_cell[    3024] = 32'h00000000;
        ram_cell[    3025] = 32'h00000000;
        ram_cell[    3026] = 32'h00000000;
        ram_cell[    3027] = 32'h00000000;
        ram_cell[    3028] = 32'h00000000;
        ram_cell[    3029] = 32'h00000000;
        ram_cell[    3030] = 32'h00000000;
        ram_cell[    3031] = 32'h00000000;
        ram_cell[    3032] = 32'h00000000;
        ram_cell[    3033] = 32'h00000000;
        ram_cell[    3034] = 32'h00000000;
        ram_cell[    3035] = 32'h00000000;
        ram_cell[    3036] = 32'h00000000;
        ram_cell[    3037] = 32'h00000000;
        ram_cell[    3038] = 32'h00000000;
        ram_cell[    3039] = 32'h00000000;
        ram_cell[    3040] = 32'h00000000;
        ram_cell[    3041] = 32'h00000000;
        ram_cell[    3042] = 32'h00000000;
        ram_cell[    3043] = 32'h00000000;
        ram_cell[    3044] = 32'h00000000;
        ram_cell[    3045] = 32'h00000000;
        ram_cell[    3046] = 32'h00000000;
        ram_cell[    3047] = 32'h00000000;
        ram_cell[    3048] = 32'h00000000;
        ram_cell[    3049] = 32'h00000000;
        ram_cell[    3050] = 32'h00000000;
        ram_cell[    3051] = 32'h00000000;
        ram_cell[    3052] = 32'h00000000;
        ram_cell[    3053] = 32'h00000000;
        ram_cell[    3054] = 32'h00000000;
        ram_cell[    3055] = 32'h00000000;
        ram_cell[    3056] = 32'h00000000;
        ram_cell[    3057] = 32'h00000000;
        ram_cell[    3058] = 32'h00000000;
        ram_cell[    3059] = 32'h00000000;
        ram_cell[    3060] = 32'h00000000;
        ram_cell[    3061] = 32'h00000000;
        ram_cell[    3062] = 32'h00000000;
        ram_cell[    3063] = 32'h00000000;
        ram_cell[    3064] = 32'h00000000;
        ram_cell[    3065] = 32'h00000000;
        ram_cell[    3066] = 32'h00000000;
        ram_cell[    3067] = 32'h00000000;
        ram_cell[    3068] = 32'h00000000;
        ram_cell[    3069] = 32'h00000000;
        ram_cell[    3070] = 32'h00000000;
        ram_cell[    3071] = 32'h00000000;
        ram_cell[    3072] = 32'h00000000;
        ram_cell[    3073] = 32'h00000000;
        ram_cell[    3074] = 32'h00000000;
        ram_cell[    3075] = 32'h00000000;
        ram_cell[    3076] = 32'h00000000;
        ram_cell[    3077] = 32'h00000000;
        ram_cell[    3078] = 32'h00000000;
        ram_cell[    3079] = 32'h00000000;
        ram_cell[    3080] = 32'h00000000;
        ram_cell[    3081] = 32'h00000000;
        ram_cell[    3082] = 32'h00000000;
        ram_cell[    3083] = 32'h00000000;
        ram_cell[    3084] = 32'h00000000;
        ram_cell[    3085] = 32'h00000000;
        ram_cell[    3086] = 32'h00000000;
        ram_cell[    3087] = 32'h00000000;
        ram_cell[    3088] = 32'h00000000;
        ram_cell[    3089] = 32'h00000000;
        ram_cell[    3090] = 32'h00000000;
        ram_cell[    3091] = 32'h00000000;
        ram_cell[    3092] = 32'h00000000;
        ram_cell[    3093] = 32'h00000000;
        ram_cell[    3094] = 32'h00000000;
        ram_cell[    3095] = 32'h00000000;
        ram_cell[    3096] = 32'h00000000;
        ram_cell[    3097] = 32'h00000000;
        ram_cell[    3098] = 32'h00000000;
        ram_cell[    3099] = 32'h00000000;
        ram_cell[    3100] = 32'h00000000;
        ram_cell[    3101] = 32'h00000000;
        ram_cell[    3102] = 32'h00000000;
        ram_cell[    3103] = 32'h00000000;
        ram_cell[    3104] = 32'h00000000;
        ram_cell[    3105] = 32'h00000000;
        ram_cell[    3106] = 32'h00000000;
        ram_cell[    3107] = 32'h00000000;
        ram_cell[    3108] = 32'h00000000;
        ram_cell[    3109] = 32'h00000000;
        ram_cell[    3110] = 32'h00000000;
        ram_cell[    3111] = 32'h00000000;
        ram_cell[    3112] = 32'h00000000;
        ram_cell[    3113] = 32'h00000000;
        ram_cell[    3114] = 32'h00000000;
        ram_cell[    3115] = 32'h00000000;
        ram_cell[    3116] = 32'h00000000;
        ram_cell[    3117] = 32'h00000000;
        ram_cell[    3118] = 32'h00000000;
        ram_cell[    3119] = 32'h00000000;
        ram_cell[    3120] = 32'h00000000;
        ram_cell[    3121] = 32'h00000000;
        ram_cell[    3122] = 32'h00000000;
        ram_cell[    3123] = 32'h00000000;
        ram_cell[    3124] = 32'h00000000;
        ram_cell[    3125] = 32'h00000000;
        ram_cell[    3126] = 32'h00000000;
        ram_cell[    3127] = 32'h00000000;
        ram_cell[    3128] = 32'h00000000;
        ram_cell[    3129] = 32'h00000000;
        ram_cell[    3130] = 32'h00000000;
        ram_cell[    3131] = 32'h00000000;
        ram_cell[    3132] = 32'h00000000;
        ram_cell[    3133] = 32'h00000000;
        ram_cell[    3134] = 32'h00000000;
        ram_cell[    3135] = 32'h00000000;
        ram_cell[    3136] = 32'h00000000;
        ram_cell[    3137] = 32'h00000000;
        ram_cell[    3138] = 32'h00000000;
        ram_cell[    3139] = 32'h00000000;
        ram_cell[    3140] = 32'h00000000;
        ram_cell[    3141] = 32'h00000000;
        ram_cell[    3142] = 32'h00000000;
        ram_cell[    3143] = 32'h00000000;
        ram_cell[    3144] = 32'h00000000;
        ram_cell[    3145] = 32'h00000000;
        ram_cell[    3146] = 32'h00000000;
        ram_cell[    3147] = 32'h00000000;
        ram_cell[    3148] = 32'h00000000;
        ram_cell[    3149] = 32'h00000000;
        ram_cell[    3150] = 32'h00000000;
        ram_cell[    3151] = 32'h00000000;
        ram_cell[    3152] = 32'h00000000;
        ram_cell[    3153] = 32'h00000000;
        ram_cell[    3154] = 32'h00000000;
        ram_cell[    3155] = 32'h00000000;
        ram_cell[    3156] = 32'h00000000;
        ram_cell[    3157] = 32'h00000000;
        ram_cell[    3158] = 32'h00000000;
        ram_cell[    3159] = 32'h00000000;
        ram_cell[    3160] = 32'h00000000;
        ram_cell[    3161] = 32'h00000000;
        ram_cell[    3162] = 32'h00000000;
        ram_cell[    3163] = 32'h00000000;
        ram_cell[    3164] = 32'h00000000;
        ram_cell[    3165] = 32'h00000000;
        ram_cell[    3166] = 32'h00000000;
        ram_cell[    3167] = 32'h00000000;
        ram_cell[    3168] = 32'h00000000;
        ram_cell[    3169] = 32'h00000000;
        ram_cell[    3170] = 32'h00000000;
        ram_cell[    3171] = 32'h00000000;
        ram_cell[    3172] = 32'h00000000;
        ram_cell[    3173] = 32'h00000000;
        ram_cell[    3174] = 32'h00000000;
        ram_cell[    3175] = 32'h00000000;
        ram_cell[    3176] = 32'h00000000;
        ram_cell[    3177] = 32'h00000000;
        ram_cell[    3178] = 32'h00000000;
        ram_cell[    3179] = 32'h00000000;
        ram_cell[    3180] = 32'h00000000;
        ram_cell[    3181] = 32'h00000000;
        ram_cell[    3182] = 32'h00000000;
        ram_cell[    3183] = 32'h00000000;
        ram_cell[    3184] = 32'h00000000;
        ram_cell[    3185] = 32'h00000000;
        ram_cell[    3186] = 32'h00000000;
        ram_cell[    3187] = 32'h00000000;
        ram_cell[    3188] = 32'h00000000;
        ram_cell[    3189] = 32'h00000000;
        ram_cell[    3190] = 32'h00000000;
        ram_cell[    3191] = 32'h00000000;
        ram_cell[    3192] = 32'h00000000;
        ram_cell[    3193] = 32'h00000000;
        ram_cell[    3194] = 32'h00000000;
        ram_cell[    3195] = 32'h00000000;
        ram_cell[    3196] = 32'h00000000;
        ram_cell[    3197] = 32'h00000000;
        ram_cell[    3198] = 32'h00000000;
        ram_cell[    3199] = 32'h00000000;
        ram_cell[    3200] = 32'h00000000;
        ram_cell[    3201] = 32'h00000000;
        ram_cell[    3202] = 32'h00000000;
        ram_cell[    3203] = 32'h00000000;
        ram_cell[    3204] = 32'h00000000;
        ram_cell[    3205] = 32'h00000000;
        ram_cell[    3206] = 32'h00000000;
        ram_cell[    3207] = 32'h00000000;
        ram_cell[    3208] = 32'h00000000;
        ram_cell[    3209] = 32'h00000000;
        ram_cell[    3210] = 32'h00000000;
        ram_cell[    3211] = 32'h00000000;
        ram_cell[    3212] = 32'h00000000;
        ram_cell[    3213] = 32'h00000000;
        ram_cell[    3214] = 32'h00000000;
        ram_cell[    3215] = 32'h00000000;
        ram_cell[    3216] = 32'h00000000;
        ram_cell[    3217] = 32'h00000000;
        ram_cell[    3218] = 32'h00000000;
        ram_cell[    3219] = 32'h00000000;
        ram_cell[    3220] = 32'h00000000;
        ram_cell[    3221] = 32'h00000000;
        ram_cell[    3222] = 32'h00000000;
        ram_cell[    3223] = 32'h00000000;
        ram_cell[    3224] = 32'h00000000;
        ram_cell[    3225] = 32'h00000000;
        ram_cell[    3226] = 32'h00000000;
        ram_cell[    3227] = 32'h00000000;
        ram_cell[    3228] = 32'h00000000;
        ram_cell[    3229] = 32'h00000000;
        ram_cell[    3230] = 32'h00000000;
        ram_cell[    3231] = 32'h00000000;
        ram_cell[    3232] = 32'h00000000;
        ram_cell[    3233] = 32'h00000000;
        ram_cell[    3234] = 32'h00000000;
        ram_cell[    3235] = 32'h00000000;
        ram_cell[    3236] = 32'h00000000;
        ram_cell[    3237] = 32'h00000000;
        ram_cell[    3238] = 32'h00000000;
        ram_cell[    3239] = 32'h00000000;
        ram_cell[    3240] = 32'h00000000;
        ram_cell[    3241] = 32'h00000000;
        ram_cell[    3242] = 32'h00000000;
        ram_cell[    3243] = 32'h00000000;
        ram_cell[    3244] = 32'h00000000;
        ram_cell[    3245] = 32'h00000000;
        ram_cell[    3246] = 32'h00000000;
        ram_cell[    3247] = 32'h00000000;
        ram_cell[    3248] = 32'h00000000;
        ram_cell[    3249] = 32'h00000000;
        ram_cell[    3250] = 32'h00000000;
        ram_cell[    3251] = 32'h00000000;
        ram_cell[    3252] = 32'h00000000;
        ram_cell[    3253] = 32'h00000000;
        ram_cell[    3254] = 32'h00000000;
        ram_cell[    3255] = 32'h00000000;
        ram_cell[    3256] = 32'h00000000;
        ram_cell[    3257] = 32'h00000000;
        ram_cell[    3258] = 32'h00000000;
        ram_cell[    3259] = 32'h00000000;
        ram_cell[    3260] = 32'h00000000;
        ram_cell[    3261] = 32'h00000000;
        ram_cell[    3262] = 32'h00000000;
        ram_cell[    3263] = 32'h00000000;
        ram_cell[    3264] = 32'h00000000;
        ram_cell[    3265] = 32'h00000000;
        ram_cell[    3266] = 32'h00000000;
        ram_cell[    3267] = 32'h00000000;
        ram_cell[    3268] = 32'h0ff000ff;
        ram_cell[    3269] = 32'hefefefef;
        ram_cell[    3270] = 32'hefefefef;
        ram_cell[    3271] = 32'h0000efef;
        ram_cell[    3272] = 32'hff0000ff;
        ram_cell[    3273] = 32'hf00f0ff0;
        ram_cell[    3274] = 32'hbeefbeef;
        ram_cell[    3275] = 32'hbeefbeef;
        ram_cell[    3276] = 32'hbeefbeef;
        ram_cell[    3277] = 32'hbeefbeef;
        ram_cell[    3278] = 32'hbeefbeef;
        ram_cell[    3279] = 32'h00000000;
        ram_cell[    3280] = 32'h00ff00ff;
        ram_cell[    3281] = 32'hff00ff00;
        ram_cell[    3282] = 32'h0ff00ff0;
        ram_cell[    3283] = 32'hf00ff00f;
        ram_cell[    3284] = 32'hdeadbeef;
        ram_cell[    3285] = 32'hdeadbeef;
        ram_cell[    3286] = 32'hdeadbeef;
        ram_cell[    3287] = 32'hdeadbeef;
        ram_cell[    3288] = 32'hdeadbeef;
        ram_cell[    3289] = 32'hdeadbeef;
        ram_cell[    3290] = 32'hdeadbeef;
        ram_cell[    3291] = 32'hdeadbeef;
        ram_cell[    3292] = 32'hdeadbeef;
        ram_cell[    3293] = 32'hdeadbeef;
        ram_cell[    3294] = 32'h00000000;
        ram_cell[    3295] = 32'h00000000;
        ram_cell[    3296] = 32'h14d68693;
        ram_cell[    3297] = 32'h00000000;
        ram_cell[    3298] = 32'h00000000;
        ram_cell[    3299] = 32'h00000000;
        ram_cell[    3300] = 32'h00000000;
        ram_cell[    3301] = 32'h00000000;
        ram_cell[    3302] = 32'h00000000;
        ram_cell[    3303] = 32'h00000000;
        ram_cell[    3304] = 32'h00000000;
        ram_cell[    3305] = 32'h00000000;
        ram_cell[    3306] = 32'h00000000;
        ram_cell[    3307] = 32'h00000000;
        ram_cell[    3308] = 32'h00000000;
        ram_cell[    3309] = 32'h00000000;
        ram_cell[    3310] = 32'h00000000;
        ram_cell[    3311] = 32'h00000000;
        ram_cell[    3312] = 32'h00000000;
        ram_cell[    3313] = 32'h00000000;
        ram_cell[    3314] = 32'h00000000;
        ram_cell[    3315] = 32'h00000000;
        ram_cell[    3316] = 32'h00000000;
        ram_cell[    3317] = 32'h00000000;
        ram_cell[    3318] = 32'h00000000;
        ram_cell[    3319] = 32'h00000000;
        ram_cell[    3320] = 32'h00000000;
        ram_cell[    3321] = 32'h00000000;
        ram_cell[    3322] = 32'h00000000;
        ram_cell[    3323] = 32'h00000000;
        ram_cell[    3324] = 32'h00000000;
        ram_cell[    3325] = 32'h00000000;
        ram_cell[    3326] = 32'h00000000;
        ram_cell[    3327] = 32'h00000000;
        ram_cell[    3328] = 32'h00000000;
        ram_cell[    3329] = 32'h00000000;
end

endmodule
